//Generate the verilog at 2024-03-17T16:07:49
module top (
clk,
ps2_clk,
ps2_data,
rst_n,
ascii_code,
data,
value_seg
);

input clk ;
input ps2_clk ;
input ps2_data ;
input rst_n ;
output [7:0] ascii_code ;
output [7:0] data ;
output [41:0] value_seg ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire _143_ ;
wire _144_ ;
wire _145_ ;
wire _146_ ;
wire _147_ ;
wire _148_ ;
wire _149_ ;
wire _150_ ;
wire _151_ ;
wire _152_ ;
wire _153_ ;
wire _154_ ;
wire _155_ ;
wire _156_ ;
wire _157_ ;
wire _158_ ;
wire _159_ ;
wire _160_ ;
wire _161_ ;
wire _162_ ;
wire _163_ ;
wire _164_ ;
wire _165_ ;
wire _166_ ;
wire _167_ ;
wire _168_ ;
wire _169_ ;
wire _170_ ;
wire _171_ ;
wire _172_ ;
wire _173_ ;
wire _174_ ;
wire _175_ ;
wire _176_ ;
wire _177_ ;
wire _178_ ;
wire _179_ ;
wire _180_ ;
wire _181_ ;
wire _182_ ;
wire _183_ ;
wire _184_ ;
wire _185_ ;
wire _186_ ;
wire _187_ ;
wire _188_ ;
wire _189_ ;
wire _190_ ;
wire _191_ ;
wire _192_ ;
wire _193_ ;
wire _194_ ;
wire _195_ ;
wire _196_ ;
wire _197_ ;
wire _198_ ;
wire _199_ ;
wire _200_ ;
wire _201_ ;
wire _202_ ;
wire _203_ ;
wire _204_ ;
wire _205_ ;
wire _206_ ;
wire _207_ ;
wire _208_ ;
wire _209_ ;
wire _210_ ;
wire _211_ ;
wire _212_ ;
wire _213_ ;
wire _214_ ;
wire _215_ ;
wire _216_ ;
wire _217_ ;
wire _218_ ;
wire _219_ ;
wire _220_ ;
wire _221_ ;
wire _222_ ;
wire _223_ ;
wire _224_ ;
wire _225_ ;
wire _226_ ;
wire _227_ ;
wire _228_ ;
wire _229_ ;
wire _230_ ;
wire _231_ ;
wire _232_ ;
wire _233_ ;
wire _234_ ;
wire _235_ ;
wire _236_ ;
wire _237_ ;
wire _238_ ;
wire _239_ ;
wire _240_ ;
wire _241_ ;
wire _242_ ;
wire _243_ ;
wire _244_ ;
wire _245_ ;
wire _246_ ;
wire _247_ ;
wire _248_ ;
wire _249_ ;
wire _250_ ;
wire _251_ ;
wire _252_ ;
wire _253_ ;
wire _254_ ;
wire _255_ ;
wire _256_ ;
wire _257_ ;
wire _258_ ;
wire _259_ ;
wire _260_ ;
wire _261_ ;
wire _262_ ;
wire _263_ ;
wire _264_ ;
wire _265_ ;
wire _266_ ;
wire _267_ ;
wire _268_ ;
wire _269_ ;
wire _270_ ;
wire _271_ ;
wire _272_ ;
wire _273_ ;
wire _274_ ;
wire _275_ ;
wire _276_ ;
wire _277_ ;
wire _278_ ;
wire _279_ ;
wire _280_ ;
wire _281_ ;
wire _282_ ;
wire _283_ ;
wire _284_ ;
wire _285_ ;
wire _286_ ;
wire _287_ ;
wire _288_ ;
wire _289_ ;
wire _290_ ;
wire _291_ ;
wire _292_ ;
wire _293_ ;
wire _294_ ;
wire _295_ ;
wire _296_ ;
wire _297_ ;
wire \buff[0] ;
wire \buff[1] ;
wire \buff[2] ;
wire \buff[3] ;
wire \buff[4] ;
wire \buff[5] ;
wire \buff[6] ;
wire \buff[7] ;
wire \count[0] ;
wire \count[1] ;
wire \count[2] ;
wire \count[3] ;
wire \count[4] ;
wire \count[5] ;
wire \count[6] ;
wire \count[7] ;
wire flag ;
wire flag_temp ;
wire \ps2_value[0] ;
wire \ps2_value[10] ;
wire \ps2_value[11] ;
wire \ps2_value[12] ;
wire \ps2_value[13] ;
wire \ps2_value[14] ;
wire \ps2_value[15] ;
wire \ps2_value[1] ;
wire \ps2_value[2] ;
wire \ps2_value[3] ;
wire \ps2_value[4] ;
wire \ps2_value[5] ;
wire \ps2_value[6] ;
wire \ps2_value[7] ;
wire \ps2_value[8] ;
wire \ps2_value[9] ;
wire \state[0] ;
wire \state[1] ;
wire \state[2] ;
wire rst_n ;
wire \data[0] ;
wire \data[1] ;
wire \data[2] ;
wire \data[3] ;
wire \data[4] ;
wire \data[5] ;
wire \data[6] ;
wire \data[7] ;
wire \ascii_code[0] ;
wire \ascii_code[1] ;
wire \ascii_code[2] ;
wire \ascii_code[3] ;
wire \ascii_code[4] ;
wire \ascii_code[5] ;
wire \ascii_code[6] ;
wire \ascii_code[7] ;
wire clk ;
wire \ScanCodeToASCII_init/_0_ ;
wire \ps2_keyboard_init/_000_ ;
wire \ps2_keyboard_init/_001_ ;
wire \ps2_keyboard_init/_002_ ;
wire \ps2_keyboard_init/_003_ ;
wire \ps2_keyboard_init/_004_ ;
wire \ps2_keyboard_init/_005_ ;
wire \ps2_keyboard_init/_006_ ;
wire \ps2_keyboard_init/_007_ ;
wire \ps2_keyboard_init/_008_ ;
wire \ps2_keyboard_init/_009_ ;
wire \ps2_keyboard_init/_010_ ;
wire \ps2_keyboard_init/_011_ ;
wire \ps2_keyboard_init/_012_ ;
wire \ps2_keyboard_init/_013_ ;
wire \ps2_keyboard_init/_014_ ;
wire \ps2_keyboard_init/_015_ ;
wire \ps2_keyboard_init/_016_ ;
wire \ps2_keyboard_init/_017_ ;
wire \ps2_keyboard_init/_018_ ;
wire \ps2_keyboard_init/_019_ ;
wire \ps2_keyboard_init/_020_ ;
wire \ps2_keyboard_init/_021_ ;
wire \ps2_keyboard_init/_022_ ;
wire \ps2_keyboard_init/_023_ ;
wire \ps2_keyboard_init/_024_ ;
wire \ps2_keyboard_init/_025_ ;
wire \ps2_keyboard_init/_026_ ;
wire \ps2_keyboard_init/_027_ ;
wire \ps2_keyboard_init/_028_ ;
wire \ps2_keyboard_init/_029_ ;
wire \ps2_keyboard_init/_030_ ;
wire \ps2_keyboard_init/_031_ ;
wire \ps2_keyboard_init/_032_ ;
wire \ps2_keyboard_init/_033_ ;
wire \ps2_keyboard_init/_034_ ;
wire \ps2_keyboard_init/_035_ ;
wire \ps2_keyboard_init/_036_ ;
wire \ps2_keyboard_init/_037_ ;
wire \ps2_keyboard_init/_038_ ;
wire \ps2_keyboard_init/_039_ ;
wire \ps2_keyboard_init/_040_ ;
wire \ps2_keyboard_init/_041_ ;
wire \ps2_keyboard_init/_042_ ;
wire \ps2_keyboard_init/_043_ ;
wire \ps2_keyboard_init/_044_ ;
wire \ps2_keyboard_init/_045_ ;
wire \ps2_keyboard_init/_046_ ;
wire \ps2_keyboard_init/_047_ ;
wire \ps2_keyboard_init/_048_ ;
wire \ps2_keyboard_init/_049_ ;
wire \ps2_keyboard_init/_050_ ;
wire \ps2_keyboard_init/_051_ ;
wire \ps2_keyboard_init/_052_ ;
wire \ps2_keyboard_init/_053_ ;
wire \ps2_keyboard_init/_054_ ;
wire \ps2_keyboard_init/_055_ ;
wire \ps2_keyboard_init/_056_ ;
wire \ps2_keyboard_init/_057_ ;
wire \ps2_keyboard_init/_058_ ;
wire \ps2_keyboard_init/_059_ ;
wire \ps2_keyboard_init/_060_ ;
wire \ps2_keyboard_init/_061_ ;
wire \ps2_keyboard_init/_062_ ;
wire \ps2_keyboard_init/_063_ ;
wire \ps2_keyboard_init/_064_ ;
wire \ps2_keyboard_init/_065_ ;
wire \ps2_keyboard_init/_066_ ;
wire \ps2_keyboard_init/_067_ ;
wire \ps2_keyboard_init/_068_ ;
wire \ps2_keyboard_init/_069_ ;
wire \ps2_keyboard_init/_070_ ;
wire \ps2_keyboard_init/_071_ ;
wire \ps2_keyboard_init/_072_ ;
wire \ps2_keyboard_init/_073_ ;
wire \ps2_keyboard_init/_074_ ;
wire \ps2_keyboard_init/_075_ ;
wire \ps2_keyboard_init/_076_ ;
wire \ps2_keyboard_init/_077_ ;
wire \ps2_keyboard_init/_078_ ;
wire \ps2_keyboard_init/_079_ ;
wire \ps2_keyboard_init/_080_ ;
wire \ps2_keyboard_init/_081_ ;
wire \ps2_keyboard_init/_082_ ;
wire \ps2_keyboard_init/_083_ ;
wire \ps2_keyboard_init/_084_ ;
wire \ps2_keyboard_init/_085_ ;
wire \ps2_keyboard_init/_086_ ;
wire \ps2_keyboard_init/_087_ ;
wire \ps2_keyboard_init/_088_ ;
wire \ps2_keyboard_init/_089_ ;
wire \ps2_keyboard_init/_090_ ;
wire \ps2_keyboard_init/_091_ ;
wire \ps2_keyboard_init/_092_ ;
wire \ps2_keyboard_init/_093_ ;
wire \ps2_keyboard_init/_094_ ;
wire \ps2_keyboard_init/_095_ ;
wire \ps2_keyboard_init/_096_ ;
wire \ps2_keyboard_init/_097_ ;
wire \ps2_keyboard_init/_098_ ;
wire \ps2_keyboard_init/_099_ ;
wire \ps2_keyboard_init/_100_ ;
wire \ps2_keyboard_init/_101_ ;
wire \ps2_keyboard_init/_102_ ;
wire \ps2_keyboard_init/_103_ ;
wire \ps2_keyboard_init/_104_ ;
wire \ps2_keyboard_init/_105_ ;
wire \ps2_keyboard_init/_106_ ;
wire \ps2_keyboard_init/_107_ ;
wire \ps2_keyboard_init/_108_ ;
wire \ps2_keyboard_init/_109_ ;
wire \ps2_keyboard_init/_110_ ;
wire \ps2_keyboard_init/_111_ ;
wire \ps2_keyboard_init/_112_ ;
wire \ps2_keyboard_init/_113_ ;
wire \ps2_keyboard_init/_114_ ;
wire \ps2_keyboard_init/_115_ ;
wire \ps2_keyboard_init/_116_ ;
wire \ps2_keyboard_init/_117_ ;
wire \ps2_keyboard_init/_118_ ;
wire \ps2_keyboard_init/_119_ ;
wire \ps2_keyboard_init/_120_ ;
wire \ps2_keyboard_init/_121_ ;
wire \ps2_keyboard_init/_122_ ;
wire \ps2_keyboard_init/_123_ ;
wire \ps2_keyboard_init/_124_ ;
wire \ps2_keyboard_init/_125_ ;
wire \ps2_keyboard_init/_126_ ;
wire \ps2_keyboard_init/_127_ ;
wire \ps2_keyboard_init/_128_ ;
wire \ps2_keyboard_init/_129_ ;
wire \ps2_keyboard_init/_130_ ;
wire \ps2_keyboard_init/_131_ ;
wire \ps2_keyboard_init/_132_ ;
wire \ps2_keyboard_init/_133_ ;
wire \ps2_keyboard_init/_134_ ;
wire \ps2_keyboard_init/_135_ ;
wire \ps2_keyboard_init/_136_ ;
wire \ps2_keyboard_init/_137_ ;
wire \ps2_keyboard_init/_138_ ;
wire \ps2_keyboard_init/_139_ ;
wire \ps2_keyboard_init/_140_ ;
wire \ps2_keyboard_init/_141_ ;
wire \ps2_keyboard_init/_142_ ;
wire \ps2_keyboard_init/_143_ ;
wire \ps2_keyboard_init/_144_ ;
wire \ps2_keyboard_init/_145_ ;
wire \ps2_keyboard_init/_146_ ;
wire \ps2_keyboard_init/_147_ ;
wire \ps2_keyboard_init/_148_ ;
wire \ps2_keyboard_init/_149_ ;
wire \ps2_keyboard_init/_150_ ;
wire \ps2_keyboard_init/_151_ ;
wire \ps2_keyboard_init/_152_ ;
wire \ps2_keyboard_init/_153_ ;
wire \ps2_keyboard_init/_154_ ;
wire \ps2_keyboard_init/_155_ ;
wire \ps2_keyboard_init/_156_ ;
wire \ps2_keyboard_init/_157_ ;
wire \ps2_keyboard_init/_158_ ;
wire \ps2_keyboard_init/_159_ ;
wire \ps2_keyboard_init/_160_ ;
wire \ps2_keyboard_init/_161_ ;
wire \ps2_keyboard_init/_162_ ;
wire \ps2_keyboard_init/_163_ ;
wire \ps2_keyboard_init/_164_ ;
wire \ps2_keyboard_init/_165_ ;
wire \ps2_keyboard_init/_166_ ;
wire \ps2_keyboard_init/_167_ ;
wire \ps2_keyboard_init/_168_ ;
wire \ps2_keyboard_init/_169_ ;
wire \ps2_keyboard_init/_170_ ;
wire \ps2_keyboard_init/_171_ ;
wire \ps2_keyboard_init/buffer[0] ;
wire \ps2_keyboard_init/buffer[1] ;
wire \ps2_keyboard_init/buffer[2] ;
wire \ps2_keyboard_init/buffer[3] ;
wire \ps2_keyboard_init/buffer[4] ;
wire \ps2_keyboard_init/buffer[5] ;
wire \ps2_keyboard_init/buffer[6] ;
wire \ps2_keyboard_init/buffer[7] ;
wire \ps2_keyboard_init/buffer[8] ;
wire \ps2_keyboard_init/buffer[9] ;
wire \ps2_keyboard_init/count[0] ;
wire \ps2_keyboard_init/count[1] ;
wire \ps2_keyboard_init/count[2] ;
wire \ps2_keyboard_init/count[3] ;
wire \ps2_keyboard_init/ps2_clk_sync[0] ;
wire \ps2_keyboard_init/ps2_clk_sync[1] ;
wire \ps2_keyboard_init/ps2_clk_sync[2] ;
wire ps2_data ;
wire ps2_clk ;
wire \seg0/_00_ ;
wire \seg0/_01_ ;
wire \seg0/_02_ ;
wire \seg0/_03_ ;
wire \seg0/_04_ ;
wire \seg0/_05_ ;
wire \seg0/_06_ ;
wire \seg0/_07_ ;
wire \seg0/_08_ ;
wire \seg0/_09_ ;
wire \seg0/_10_ ;
wire \seg0/_11_ ;
wire \seg0/_12_ ;
wire \seg0/_13_ ;
wire \seg0/_14_ ;
wire \seg0/_15_ ;
wire \seg0/_16_ ;
wire \seg0/_17_ ;
wire \seg0/_18_ ;
wire \seg0/_19_ ;
wire \seg0/_20_ ;
wire \seg0/_21_ ;
wire \seg0/_22_ ;
wire \seg0/_23_ ;
wire \seg0/_24_ ;
wire \seg0/_25_ ;
wire \seg0/_26_ ;
wire \seg0/_27_ ;
wire \seg0/_28_ ;
wire \seg0/_29_ ;
wire \seg0/_30_ ;
wire \seg0/_31_ ;
wire \seg0/_32_ ;
wire \seg0/_33_ ;
wire \seg0/_34_ ;
wire \seg0/_35_ ;
wire \seg0/_36_ ;
wire \seg0/_37_ ;
wire \value_seg[0] ;
wire \value_seg[1] ;
wire \value_seg[2] ;
wire \value_seg[3] ;
wire \value_seg[4] ;
wire \value_seg[5] ;
wire \value_seg[6] ;
wire \seg1/_00_ ;
wire \seg1/_01_ ;
wire \seg1/_02_ ;
wire \seg1/_03_ ;
wire \seg1/_04_ ;
wire \seg1/_05_ ;
wire \seg1/_06_ ;
wire \seg1/_07_ ;
wire \seg1/_08_ ;
wire \seg1/_09_ ;
wire \seg1/_10_ ;
wire \seg1/_11_ ;
wire \seg1/_12_ ;
wire \seg1/_13_ ;
wire \seg1/_14_ ;
wire \seg1/_15_ ;
wire \seg1/_16_ ;
wire \seg1/_17_ ;
wire \seg1/_18_ ;
wire \seg1/_19_ ;
wire \seg1/_20_ ;
wire \seg1/_21_ ;
wire \seg1/_22_ ;
wire \seg1/_23_ ;
wire \seg1/_24_ ;
wire \seg1/_25_ ;
wire \seg1/_26_ ;
wire \seg1/_27_ ;
wire \seg1/_28_ ;
wire \seg1/_29_ ;
wire \seg1/_30_ ;
wire \seg1/_31_ ;
wire \seg1/_32_ ;
wire \seg1/_33_ ;
wire \seg1/_34_ ;
wire \seg1/_35_ ;
wire \seg1/_36_ ;
wire \seg1/_37_ ;
wire \value_seg[7] ;
wire \value_seg[8] ;
wire \value_seg[9] ;
wire \value_seg[10] ;
wire \value_seg[11] ;
wire \value_seg[12] ;
wire \value_seg[13] ;
wire \seg2/_00_ ;
wire \seg2/_01_ ;
wire \seg2/_02_ ;
wire \seg2/_03_ ;
wire \seg2/_04_ ;
wire \seg2/_05_ ;
wire \seg2/_06_ ;
wire \seg2/_07_ ;
wire \seg2/_08_ ;
wire \seg2/_09_ ;
wire \seg2/_10_ ;
wire \seg2/_11_ ;
wire \seg2/_12_ ;
wire \seg2/_13_ ;
wire \seg2/_14_ ;
wire \seg2/_15_ ;
wire \seg2/_16_ ;
wire \seg2/_17_ ;
wire \seg2/_18_ ;
wire \seg2/_19_ ;
wire \seg2/_20_ ;
wire \seg2/_21_ ;
wire \seg2/_22_ ;
wire \seg2/_23_ ;
wire \seg2/_24_ ;
wire \seg2/_25_ ;
wire \seg2/_26_ ;
wire \seg2/_27_ ;
wire \seg2/_28_ ;
wire \seg2/_29_ ;
wire \seg2/_30_ ;
wire \seg2/_31_ ;
wire \seg2/_32_ ;
wire \seg2/_33_ ;
wire \seg2/_34_ ;
wire \seg2/_35_ ;
wire \seg2/_36_ ;
wire \seg2/_37_ ;
wire \value_seg[14] ;
wire \value_seg[15] ;
wire \value_seg[16] ;
wire \value_seg[17] ;
wire \value_seg[18] ;
wire \value_seg[19] ;
wire \value_seg[20] ;
wire \seg3/_00_ ;
wire \seg3/_01_ ;
wire \seg3/_02_ ;
wire \seg3/_03_ ;
wire \seg3/_04_ ;
wire \seg3/_05_ ;
wire \seg3/_06_ ;
wire \seg3/_07_ ;
wire \seg3/_08_ ;
wire \seg3/_09_ ;
wire \seg3/_10_ ;
wire \seg3/_11_ ;
wire \seg3/_12_ ;
wire \seg3/_13_ ;
wire \seg3/_14_ ;
wire \seg3/_15_ ;
wire \seg3/_16_ ;
wire \seg3/_17_ ;
wire \seg3/_18_ ;
wire \seg3/_19_ ;
wire \seg3/_20_ ;
wire \seg3/_21_ ;
wire \seg3/_22_ ;
wire \seg3/_23_ ;
wire \seg3/_24_ ;
wire \seg3/_25_ ;
wire \seg3/_26_ ;
wire \seg3/_27_ ;
wire \seg3/_28_ ;
wire \seg3/_29_ ;
wire \seg3/_30_ ;
wire \seg3/_31_ ;
wire \seg3/_32_ ;
wire \seg3/_33_ ;
wire \seg3/_34_ ;
wire \seg3/_35_ ;
wire \seg3/_36_ ;
wire \seg3/_37_ ;
wire \value_seg[21] ;
wire \value_seg[22] ;
wire \value_seg[23] ;
wire \value_seg[24] ;
wire \value_seg[25] ;
wire \value_seg[26] ;
wire \value_seg[27] ;
wire \seg4/_00_ ;
wire \seg4/_01_ ;
wire \seg4/_02_ ;
wire \seg4/_03_ ;
wire \seg4/_04_ ;
wire \seg4/_05_ ;
wire \seg4/_06_ ;
wire \seg4/_07_ ;
wire \seg4/_08_ ;
wire \seg4/_09_ ;
wire \seg4/_10_ ;
wire \seg4/_11_ ;
wire \seg4/_12_ ;
wire \seg4/_13_ ;
wire \seg4/_14_ ;
wire \seg4/_15_ ;
wire \seg4/_16_ ;
wire \seg4/_17_ ;
wire \seg4/_18_ ;
wire \seg4/_19_ ;
wire \seg4/_20_ ;
wire \seg4/_21_ ;
wire \seg4/_22_ ;
wire \seg4/_23_ ;
wire \seg4/_24_ ;
wire \seg4/_25_ ;
wire \seg4/_26_ ;
wire \seg4/_27_ ;
wire \seg4/_28_ ;
wire \seg4/_29_ ;
wire \seg4/_30_ ;
wire \seg4/_31_ ;
wire \seg4/_32_ ;
wire \seg4/_33_ ;
wire \seg4/_34_ ;
wire \seg4/_35_ ;
wire \seg4/_36_ ;
wire \seg4/_37_ ;
wire \value_seg[28] ;
wire \value_seg[29] ;
wire \value_seg[30] ;
wire \value_seg[31] ;
wire \value_seg[32] ;
wire \value_seg[33] ;
wire \value_seg[34] ;
wire \seg5/_00_ ;
wire \seg5/_01_ ;
wire \seg5/_02_ ;
wire \seg5/_03_ ;
wire \seg5/_04_ ;
wire \seg5/_05_ ;
wire \seg5/_06_ ;
wire \seg5/_07_ ;
wire \seg5/_08_ ;
wire \seg5/_09_ ;
wire \seg5/_10_ ;
wire \seg5/_11_ ;
wire \seg5/_12_ ;
wire \seg5/_13_ ;
wire \seg5/_14_ ;
wire \seg5/_15_ ;
wire \seg5/_16_ ;
wire \seg5/_17_ ;
wire \seg5/_18_ ;
wire \seg5/_19_ ;
wire \seg5/_20_ ;
wire \seg5/_21_ ;
wire \seg5/_22_ ;
wire \seg5/_23_ ;
wire \seg5/_24_ ;
wire \seg5/_25_ ;
wire \seg5/_26_ ;
wire \seg5/_27_ ;
wire \seg5/_28_ ;
wire \seg5/_29_ ;
wire \seg5/_30_ ;
wire \seg5/_31_ ;
wire \seg5/_32_ ;
wire \seg5/_33_ ;
wire \seg5/_34_ ;
wire \seg5/_35_ ;
wire \seg5/_36_ ;
wire \seg5/_37_ ;
wire \value_seg[35] ;
wire \value_seg[36] ;
wire \value_seg[37] ;
wire \value_seg[38] ;
wire \value_seg[39] ;
wire \value_seg[40] ;
wire \value_seg[41] ;

XNOR2_X1 _298_ ( .A(_125_ ), .B(_140_ ), .ZN(_143_ ) );
XNOR2_X1 _299_ ( .A(_124_ ), .B(_139_ ), .ZN(_144_ ) );
XNOR2_X1 _300_ ( .A(_121_ ), .B(_136_ ), .ZN(_145_ ) );
XNOR2_X1 _301_ ( .A(_120_ ), .B(_135_ ), .ZN(_146_ ) );
AND4_X1 _302_ ( .A1(_143_ ), .A2(_144_ ), .A3(_145_ ), .A4(_146_ ), .ZN(_147_ ) );
XNOR2_X1 _303_ ( .A(_122_ ), .B(_137_ ), .ZN(_148_ ) );
XNOR2_X1 _304_ ( .A(_118_ ), .B(_133_ ), .ZN(_149_ ) );
XNOR2_X1 _305_ ( .A(_123_ ), .B(_138_ ), .ZN(_150_ ) );
XNOR2_X1 _306_ ( .A(_119_ ), .B(_134_ ), .ZN(_151_ ) );
AND4_X1 _307_ ( .A1(_148_ ), .A2(_149_ ), .A3(_150_ ), .A4(_151_ ), .ZN(_152_ ) );
INV_X1 _308_ ( .A(_277_ ), .ZN(_153_ ) );
NAND3_X1 _309_ ( .A1(_147_ ), .A2(_152_ ), .A3(_153_ ), .ZN(_154_ ) );
XNOR2_X1 _310_ ( .A(_142_ ), .B(_141_ ), .ZN(_155_ ) );
NAND2_X1 _311_ ( .A1(_155_ ), .A2(_153_ ), .ZN(_156_ ) );
OAI22_X1 _312_ ( .A1(_154_ ), .A2(_109_ ), .B1(_108_ ), .B2(_156_ ), .ZN(_090_ ) );
AND2_X1 _313_ ( .A1(_137_ ), .A2(_138_ ), .ZN(_157_ ) );
AND3_X4 _314_ ( .A1(_157_ ), .A2(_139_ ), .A3(_140_ ), .ZN(_158_ ) );
NOR4_X4 _315_ ( .A1(_133_ ), .A2(_134_ ), .A3(_135_ ), .A4(_136_ ), .ZN(_159_ ) );
AND2_X4 _316_ ( .A1(_158_ ), .A2(_159_ ), .ZN(_160_ ) );
OAI221_X1 _317_ ( .A(_153_ ), .B1(_108_ ), .B2(_155_ ), .C1(_160_ ), .C2(_091_ ), .ZN(_088_ ) );
AND2_X2 _318_ ( .A1(_147_ ), .A2(_152_ ), .ZN(_161_ ) );
OR3_X1 _319_ ( .A1(_161_ ), .A2(_277_ ), .A3(_109_ ), .ZN(_162_ ) );
INV_X4 _320_ ( .A(_160_ ), .ZN(_163_ ) );
OR3_X1 _321_ ( .A1(_163_ ), .A2(_277_ ), .A3(_091_ ), .ZN(_164_ ) );
NAND2_X1 _322_ ( .A1(_162_ ), .A2(_164_ ), .ZN(_089_ ) );
NAND3_X1 _323_ ( .A1(_161_ ), .A2(_153_ ), .A3(_279_ ), .ZN(_165_ ) );
MUX2_X1 _324_ ( .A(_141_ ), .B(_142_ ), .S(_165_ ), .Z(_071_ ) );
AND2_X1 _325_ ( .A1(_133_ ), .A2(_278_ ), .ZN(_166_ ) );
INV_X1 _326_ ( .A(_279_ ), .ZN(_167_ ) );
NAND2_X2 _327_ ( .A1(_167_ ), .A2(_091_ ), .ZN(_168_ ) );
NOR2_X2 _328_ ( .A1(_168_ ), .A2(_280_ ), .ZN(_169_ ) );
OR2_X2 _329_ ( .A1(_169_ ), .A2(_277_ ), .ZN(_170_ ) );
BUF_X4 _330_ ( .A(_170_ ), .Z(_171_ ) );
MUX2_X1 _331_ ( .A(_166_ ), .B(_261_ ), .S(_171_ ), .Z(_072_ ) );
AND2_X1 _332_ ( .A1(_134_ ), .A2(_278_ ), .ZN(_172_ ) );
MUX2_X1 _333_ ( .A(_172_ ), .B(_268_ ), .S(_171_ ), .Z(_079_ ) );
AND2_X1 _334_ ( .A1(_135_ ), .A2(_278_ ), .ZN(_173_ ) );
MUX2_X1 _335_ ( .A(_173_ ), .B(_269_ ), .S(_171_ ), .Z(_080_ ) );
AND2_X1 _336_ ( .A1(_136_ ), .A2(_278_ ), .ZN(_174_ ) );
MUX2_X1 _337_ ( .A(_174_ ), .B(_270_ ), .S(_171_ ), .Z(_081_ ) );
AND2_X1 _338_ ( .A1(_137_ ), .A2(_278_ ), .ZN(_175_ ) );
MUX2_X1 _339_ ( .A(_175_ ), .B(_271_ ), .S(_171_ ), .Z(_082_ ) );
AND2_X1 _340_ ( .A1(_138_ ), .A2(_278_ ), .ZN(_176_ ) );
MUX2_X1 _341_ ( .A(_176_ ), .B(_272_ ), .S(_171_ ), .Z(_083_ ) );
AND2_X1 _342_ ( .A1(_139_ ), .A2(_278_ ), .ZN(_177_ ) );
MUX2_X1 _343_ ( .A(_177_ ), .B(_273_ ), .S(_171_ ), .Z(_084_ ) );
AND2_X1 _344_ ( .A1(_140_ ), .A2(_278_ ), .ZN(_178_ ) );
MUX2_X1 _345_ ( .A(_178_ ), .B(_274_ ), .S(_171_ ), .Z(_085_ ) );
AND2_X1 _346_ ( .A1(_278_ ), .A2(_110_ ), .ZN(_179_ ) );
MUX2_X1 _347_ ( .A(_179_ ), .B(_275_ ), .S(_171_ ), .Z(_086_ ) );
AND2_X1 _348_ ( .A1(_278_ ), .A2(_111_ ), .ZN(_180_ ) );
MUX2_X1 _349_ ( .A(_180_ ), .B(_276_ ), .S(_171_ ), .Z(_087_ ) );
AND2_X1 _350_ ( .A1(_278_ ), .A2(_112_ ), .ZN(_181_ ) );
MUX2_X1 _351_ ( .A(_181_ ), .B(_262_ ), .S(_170_ ), .Z(_073_ ) );
AND2_X1 _352_ ( .A1(_278_ ), .A2(_113_ ), .ZN(_182_ ) );
MUX2_X1 _353_ ( .A(_182_ ), .B(_263_ ), .S(_170_ ), .Z(_074_ ) );
AND2_X1 _354_ ( .A1(_278_ ), .A2(_114_ ), .ZN(_183_ ) );
MUX2_X1 _355_ ( .A(_183_ ), .B(_264_ ), .S(_170_ ), .Z(_075_ ) );
AND2_X1 _356_ ( .A1(_278_ ), .A2(_115_ ), .ZN(_184_ ) );
MUX2_X1 _357_ ( .A(_184_ ), .B(_265_ ), .S(_170_ ), .Z(_076_ ) );
AND2_X1 _358_ ( .A1(_278_ ), .A2(_116_ ), .ZN(_185_ ) );
MUX2_X1 _359_ ( .A(_185_ ), .B(_266_ ), .S(_170_ ), .Z(_077_ ) );
AND2_X1 _360_ ( .A1(_278_ ), .A2(_117_ ), .ZN(_186_ ) );
MUX2_X1 _361_ ( .A(_186_ ), .B(_267_ ), .S(_170_ ), .Z(_078_ ) );
NOR3_X1 _362_ ( .A1(_168_ ), .A2(_118_ ), .A3(_280_ ), .ZN(_187_ ) );
INV_X1 _363_ ( .A(_092_ ), .ZN(_188_ ) );
NOR2_X1 _364_ ( .A1(_161_ ), .A2(_109_ ), .ZN(_189_ ) );
AND2_X4 _365_ ( .A1(_160_ ), .A2(_278_ ), .ZN(_190_ ) );
OAI21_X1 _366_ ( .A(_188_ ), .B1(_189_ ), .B2(_190_ ), .ZN(_191_ ) );
NOR2_X1 _367_ ( .A1(_155_ ), .A2(_108_ ), .ZN(_192_ ) );
AOI211_X4 _368_ ( .A(_169_ ), .B(_166_ ), .C1(_192_ ), .C2(_133_ ), .ZN(_193_ ) );
AOI211_X2 _369_ ( .A(_277_ ), .B(_187_ ), .C1(_191_ ), .C2(_193_ ), .ZN(_055_ ) );
NOR3_X1 _370_ ( .A1(_168_ ), .A2(_119_ ), .A3(_280_ ), .ZN(_194_ ) );
INV_X1 _371_ ( .A(_093_ ), .ZN(_195_ ) );
OAI21_X1 _372_ ( .A(_195_ ), .B1(_189_ ), .B2(_190_ ), .ZN(_196_ ) );
AOI211_X4 _373_ ( .A(_169_ ), .B(_172_ ), .C1(_192_ ), .C2(_134_ ), .ZN(_197_ ) );
AOI211_X2 _374_ ( .A(_277_ ), .B(_194_ ), .C1(_196_ ), .C2(_197_ ), .ZN(_056_ ) );
NOR3_X1 _375_ ( .A1(_168_ ), .A2(_120_ ), .A3(_280_ ), .ZN(_198_ ) );
INV_X1 _376_ ( .A(_094_ ), .ZN(_199_ ) );
OAI21_X1 _377_ ( .A(_199_ ), .B1(_189_ ), .B2(_190_ ), .ZN(_200_ ) );
AOI211_X4 _378_ ( .A(_169_ ), .B(_173_ ), .C1(_192_ ), .C2(_135_ ), .ZN(_201_ ) );
AOI211_X2 _379_ ( .A(_277_ ), .B(_198_ ), .C1(_200_ ), .C2(_201_ ), .ZN(_057_ ) );
NOR3_X1 _380_ ( .A1(_168_ ), .A2(_121_ ), .A3(_280_ ), .ZN(_202_ ) );
INV_X1 _381_ ( .A(_095_ ), .ZN(_203_ ) );
OAI21_X1 _382_ ( .A(_203_ ), .B1(_189_ ), .B2(_190_ ), .ZN(_204_ ) );
AOI211_X4 _383_ ( .A(_169_ ), .B(_174_ ), .C1(_192_ ), .C2(_136_ ), .ZN(_205_ ) );
AOI211_X2 _384_ ( .A(_277_ ), .B(_202_ ), .C1(_204_ ), .C2(_205_ ), .ZN(_058_ ) );
NOR3_X1 _385_ ( .A1(_168_ ), .A2(_122_ ), .A3(_280_ ), .ZN(_206_ ) );
NOR3_X1 _386_ ( .A1(_161_ ), .A2(_109_ ), .A3(_096_ ), .ZN(_207_ ) );
INV_X1 _387_ ( .A(_158_ ), .ZN(_208_ ) );
NOR3_X4 _388_ ( .A1(_208_ ), .A2(_133_ ), .A3(_136_ ), .ZN(_209_ ) );
NOR2_X1 _389_ ( .A1(_134_ ), .A2(_135_ ), .ZN(_210_ ) );
NAND3_X1 _390_ ( .A1(_209_ ), .A2(_096_ ), .A3(_210_ ), .ZN(_211_ ) );
AOI21_X1 _391_ ( .A(_207_ ), .B1(_175_ ), .B2(_211_ ), .ZN(_212_ ) );
AOI21_X1 _392_ ( .A(_169_ ), .B1(_192_ ), .B2(_137_ ), .ZN(_213_ ) );
AOI211_X4 _393_ ( .A(_277_ ), .B(_206_ ), .C1(_212_ ), .C2(_213_ ), .ZN(_059_ ) );
NOR3_X1 _394_ ( .A1(_168_ ), .A2(_123_ ), .A3(_280_ ), .ZN(_214_ ) );
NOR3_X1 _395_ ( .A1(_161_ ), .A2(_109_ ), .A3(_097_ ), .ZN(_215_ ) );
NAND3_X1 _396_ ( .A1(_209_ ), .A2(_097_ ), .A3(_210_ ), .ZN(_216_ ) );
AOI21_X1 _397_ ( .A(_215_ ), .B1(_176_ ), .B2(_216_ ), .ZN(_217_ ) );
AOI21_X1 _398_ ( .A(_169_ ), .B1(_192_ ), .B2(_138_ ), .ZN(_218_ ) );
AOI211_X4 _399_ ( .A(_277_ ), .B(_214_ ), .C1(_217_ ), .C2(_218_ ), .ZN(_060_ ) );
NOR3_X1 _400_ ( .A1(_168_ ), .A2(_124_ ), .A3(_280_ ), .ZN(_219_ ) );
NOR3_X1 _401_ ( .A1(_161_ ), .A2(_109_ ), .A3(_098_ ), .ZN(_220_ ) );
NAND3_X1 _402_ ( .A1(_209_ ), .A2(_098_ ), .A3(_210_ ), .ZN(_221_ ) );
AOI21_X1 _403_ ( .A(_220_ ), .B1(_177_ ), .B2(_221_ ), .ZN(_222_ ) );
AOI21_X1 _404_ ( .A(_169_ ), .B1(_192_ ), .B2(_139_ ), .ZN(_223_ ) );
AOI211_X4 _405_ ( .A(_277_ ), .B(_219_ ), .C1(_222_ ), .C2(_223_ ), .ZN(_061_ ) );
NOR3_X1 _406_ ( .A1(_168_ ), .A2(_125_ ), .A3(_280_ ), .ZN(_224_ ) );
NOR3_X1 _407_ ( .A1(_161_ ), .A2(_109_ ), .A3(_099_ ), .ZN(_225_ ) );
NAND3_X1 _408_ ( .A1(_209_ ), .A2(_099_ ), .A3(_210_ ), .ZN(_226_ ) );
AOI21_X1 _409_ ( .A(_225_ ), .B1(_178_ ), .B2(_226_ ), .ZN(_227_ ) );
AOI21_X1 _410_ ( .A(_169_ ), .B1(_192_ ), .B2(_140_ ), .ZN(_228_ ) );
AOI211_X4 _411_ ( .A(_277_ ), .B(_224_ ), .C1(_227_ ), .C2(_228_ ), .ZN(_062_ ) );
XNOR2_X1 _412_ ( .A(_160_ ), .B(_126_ ), .ZN(_229_ ) );
AND2_X1 _413_ ( .A1(_229_ ), .A2(_278_ ), .ZN(_230_ ) );
INV_X1 _414_ ( .A(_278_ ), .ZN(_231_ ) );
AOI211_X2 _415_ ( .A(_277_ ), .B(_230_ ), .C1(_231_ ), .C2(_100_ ), .ZN(_063_ ) );
XNOR2_X1 _416_ ( .A(_126_ ), .B(_127_ ), .ZN(_232_ ) );
AND4_X1 _417_ ( .A1(_278_ ), .A2(_209_ ), .A3(_210_ ), .A4(_232_ ), .ZN(_233_ ) );
AND2_X1 _418_ ( .A1(_209_ ), .A2(_210_ ), .ZN(_234_ ) );
AND2_X1 _419_ ( .A1(_234_ ), .A2(_278_ ), .ZN(_235_ ) );
INV_X1 _420_ ( .A(_235_ ), .ZN(_236_ ) );
AOI211_X2 _421_ ( .A(_277_ ), .B(_233_ ), .C1(_236_ ), .C2(_101_ ), .ZN(_064_ ) );
AND2_X4 _422_ ( .A1(_126_ ), .A2(_127_ ), .ZN(_237_ ) );
XNOR2_X1 _423_ ( .A(_237_ ), .B(_128_ ), .ZN(_238_ ) );
AND4_X1 _424_ ( .A1(_278_ ), .A2(_209_ ), .A3(_210_ ), .A4(_238_ ), .ZN(_239_ ) );
AOI211_X2 _425_ ( .A(_277_ ), .B(_239_ ), .C1(_236_ ), .C2(_102_ ), .ZN(_065_ ) );
AND2_X1 _426_ ( .A1(_237_ ), .A2(_128_ ), .ZN(_240_ ) );
NAND3_X1 _427_ ( .A1(_160_ ), .A2(_278_ ), .A3(_240_ ), .ZN(_241_ ) );
AND2_X1 _428_ ( .A1(_241_ ), .A2(_103_ ), .ZN(_242_ ) );
NOR2_X1 _429_ ( .A1(_241_ ), .A2(_103_ ), .ZN(_243_ ) );
NOR3_X1 _430_ ( .A1(_242_ ), .A2(_243_ ), .A3(_277_ ), .ZN(_066_ ) );
AND3_X4 _431_ ( .A1(_237_ ), .A2(_128_ ), .A3(_129_ ), .ZN(_244_ ) );
XNOR2_X1 _432_ ( .A(_244_ ), .B(_130_ ), .ZN(_245_ ) );
AND3_X1 _433_ ( .A1(_245_ ), .A2(_278_ ), .A3(_160_ ), .ZN(_246_ ) );
INV_X1 _434_ ( .A(_190_ ), .ZN(_247_ ) );
AOI211_X2 _435_ ( .A(_277_ ), .B(_246_ ), .C1(_104_ ), .C2(_247_ ), .ZN(_067_ ) );
AND2_X1 _436_ ( .A1(_244_ ), .A2(_130_ ), .ZN(_248_ ) );
INV_X1 _437_ ( .A(_248_ ), .ZN(_249_ ) );
OR4_X4 _438_ ( .A1(_231_ ), .A2(_163_ ), .A3(_249_ ), .A4(_105_ ), .ZN(_250_ ) );
NAND3_X1 _439_ ( .A1(_160_ ), .A2(_248_ ), .A3(_278_ ), .ZN(_251_ ) );
AOI21_X1 _440_ ( .A(_277_ ), .B1(_251_ ), .B2(_105_ ), .ZN(_252_ ) );
AND2_X1 _441_ ( .A1(_250_ ), .A2(_252_ ), .ZN(_068_ ) );
NAND2_X1 _442_ ( .A1(_248_ ), .A2(_131_ ), .ZN(_253_ ) );
INV_X1 _443_ ( .A(_132_ ), .ZN(_254_ ) );
NOR3_X4 _444_ ( .A1(_247_ ), .A2(_253_ ), .A3(_254_ ), .ZN(_255_ ) );
INV_X1 _445_ ( .A(_255_ ), .ZN(_256_ ) );
NAND4_X1 _446_ ( .A1(_253_ ), .A2(_278_ ), .A3(_254_ ), .A4(_160_ ), .ZN(_257_ ) );
AOI21_X1 _447_ ( .A(_277_ ), .B1(_247_ ), .B2(_106_ ), .ZN(_258_ ) );
AND3_X1 _448_ ( .A1(_256_ ), .A2(_257_ ), .A3(_258_ ), .ZN(_069_ ) );
OR2_X1 _449_ ( .A1(_255_ ), .A2(_107_ ), .ZN(_259_ ) );
NAND2_X1 _450_ ( .A1(_255_ ), .A2(_107_ ), .ZN(_260_ ) );
AOI21_X1 _451_ ( .A(_277_ ), .B1(_259_ ), .B2(_260_ ), .ZN(_070_ ) );
BUF_X1 _452_ ( .A(rst_n ), .Z(_277_ ) );
BUF_X1 _453_ ( .A(flag_temp ), .Z(_142_ ) );
BUF_X1 _454_ ( .A(flag ), .Z(_141_ ) );
BUF_X1 _455_ ( .A(\buff[0] ), .Z(_118_ ) );
BUF_X1 _456_ ( .A(\data[0] ), .Z(_133_ ) );
BUF_X1 _457_ ( .A(\buff[1] ), .Z(_119_ ) );
BUF_X1 _458_ ( .A(\data[1] ), .Z(_134_ ) );
BUF_X1 _459_ ( .A(\buff[2] ), .Z(_120_ ) );
BUF_X1 _460_ ( .A(\data[2] ), .Z(_135_ ) );
BUF_X1 _461_ ( .A(\buff[3] ), .Z(_121_ ) );
BUF_X1 _462_ ( .A(\data[3] ), .Z(_136_ ) );
BUF_X1 _463_ ( .A(\buff[4] ), .Z(_122_ ) );
BUF_X1 _464_ ( .A(\data[4] ), .Z(_137_ ) );
BUF_X1 _465_ ( .A(\buff[5] ), .Z(_123_ ) );
BUF_X1 _466_ ( .A(\data[5] ), .Z(_138_ ) );
BUF_X1 _467_ ( .A(\buff[6] ), .Z(_124_ ) );
BUF_X1 _468_ ( .A(\data[6] ), .Z(_139_ ) );
BUF_X1 _469_ ( .A(\buff[7] ), .Z(_125_ ) );
BUF_X1 _470_ ( .A(\data[7] ), .Z(_140_ ) );
BUF_X1 _471_ ( .A(_054_ ), .Z(_109_ ) );
BUF_X1 _472_ ( .A(_053_ ), .Z(_108_ ) );
BUF_X1 _473_ ( .A(_090_ ), .Z(_035_ ) );
BUF_X1 _474_ ( .A(_036_ ), .Z(_091_ ) );
BUF_X1 _475_ ( .A(_088_ ), .Z(_033_ ) );
BUF_X1 _476_ ( .A(_089_ ), .Z(_034_ ) );
BUF_X1 _477_ ( .A(\state[1] ), .Z(_279_ ) );
BUF_X1 _478_ ( .A(_071_ ), .Z(_016_ ) );
BUF_X1 _479_ ( .A(\state[2] ), .Z(_280_ ) );
BUF_X1 _480_ ( .A(\state[0] ), .Z(_278_ ) );
BUF_X1 _481_ ( .A(\ps2_value[0] ), .Z(_261_ ) );
BUF_X1 _482_ ( .A(_072_ ), .Z(_017_ ) );
BUF_X1 _483_ ( .A(\ps2_value[1] ), .Z(_268_ ) );
BUF_X1 _484_ ( .A(_079_ ), .Z(_024_ ) );
BUF_X1 _485_ ( .A(\ps2_value[2] ), .Z(_269_ ) );
BUF_X1 _486_ ( .A(_080_ ), .Z(_025_ ) );
BUF_X1 _487_ ( .A(\ps2_value[3] ), .Z(_270_ ) );
BUF_X1 _488_ ( .A(_081_ ), .Z(_026_ ) );
BUF_X1 _489_ ( .A(\ps2_value[4] ), .Z(_271_ ) );
BUF_X1 _490_ ( .A(_082_ ), .Z(_027_ ) );
BUF_X1 _491_ ( .A(\ps2_value[5] ), .Z(_272_ ) );
BUF_X1 _492_ ( .A(_083_ ), .Z(_028_ ) );
BUF_X1 _493_ ( .A(\ps2_value[6] ), .Z(_273_ ) );
BUF_X1 _494_ ( .A(_084_ ), .Z(_029_ ) );
BUF_X1 _495_ ( .A(\ps2_value[7] ), .Z(_274_ ) );
BUF_X1 _496_ ( .A(_085_ ), .Z(_030_ ) );
BUF_X1 _497_ ( .A(\ascii_code[0] ), .Z(_110_ ) );
BUF_X1 _498_ ( .A(\ps2_value[8] ), .Z(_275_ ) );
BUF_X1 _499_ ( .A(_086_ ), .Z(_031_ ) );
BUF_X1 _500_ ( .A(\ascii_code[1] ), .Z(_111_ ) );
BUF_X1 _501_ ( .A(\ps2_value[9] ), .Z(_276_ ) );
BUF_X1 _502_ ( .A(_087_ ), .Z(_032_ ) );
BUF_X1 _503_ ( .A(\ascii_code[2] ), .Z(_112_ ) );
BUF_X1 _504_ ( .A(\ps2_value[10] ), .Z(_262_ ) );
BUF_X1 _505_ ( .A(_073_ ), .Z(_018_ ) );
BUF_X1 _506_ ( .A(\ascii_code[3] ), .Z(_113_ ) );
BUF_X1 _507_ ( .A(\ps2_value[11] ), .Z(_263_ ) );
BUF_X1 _508_ ( .A(_074_ ), .Z(_019_ ) );
BUF_X1 _509_ ( .A(\ascii_code[4] ), .Z(_114_ ) );
BUF_X1 _510_ ( .A(\ps2_value[12] ), .Z(_264_ ) );
BUF_X1 _511_ ( .A(_075_ ), .Z(_020_ ) );
BUF_X1 _512_ ( .A(\ascii_code[5] ), .Z(_115_ ) );
BUF_X1 _513_ ( .A(\ps2_value[13] ), .Z(_265_ ) );
BUF_X1 _514_ ( .A(_076_ ), .Z(_021_ ) );
BUF_X1 _515_ ( .A(\ascii_code[6] ), .Z(_116_ ) );
BUF_X1 _516_ ( .A(\ps2_value[14] ), .Z(_266_ ) );
BUF_X1 _517_ ( .A(_077_ ), .Z(_022_ ) );
BUF_X1 _518_ ( .A(\ascii_code[7] ), .Z(_117_ ) );
BUF_X1 _519_ ( .A(\ps2_value[15] ), .Z(_267_ ) );
BUF_X1 _520_ ( .A(_078_ ), .Z(_023_ ) );
BUF_X1 _521_ ( .A(_037_ ), .Z(_092_ ) );
BUF_X1 _522_ ( .A(_055_ ), .Z(_000_ ) );
BUF_X1 _523_ ( .A(_038_ ), .Z(_093_ ) );
BUF_X1 _524_ ( .A(_056_ ), .Z(_001_ ) );
BUF_X1 _525_ ( .A(_039_ ), .Z(_094_ ) );
BUF_X1 _526_ ( .A(_057_ ), .Z(_002_ ) );
BUF_X1 _527_ ( .A(_040_ ), .Z(_095_ ) );
BUF_X1 _528_ ( .A(_058_ ), .Z(_003_ ) );
BUF_X1 _529_ ( .A(_041_ ), .Z(_096_ ) );
BUF_X1 _530_ ( .A(_059_ ), .Z(_004_ ) );
BUF_X1 _531_ ( .A(_042_ ), .Z(_097_ ) );
BUF_X1 _532_ ( .A(_060_ ), .Z(_005_ ) );
BUF_X1 _533_ ( .A(_043_ ), .Z(_098_ ) );
BUF_X1 _534_ ( .A(_061_ ), .Z(_006_ ) );
BUF_X1 _535_ ( .A(_044_ ), .Z(_099_ ) );
BUF_X1 _536_ ( .A(_062_ ), .Z(_007_ ) );
BUF_X1 _537_ ( .A(\count[0] ), .Z(_126_ ) );
BUF_X1 _538_ ( .A(_045_ ), .Z(_100_ ) );
BUF_X1 _539_ ( .A(_063_ ), .Z(_008_ ) );
BUF_X1 _540_ ( .A(\count[1] ), .Z(_127_ ) );
BUF_X1 _541_ ( .A(_046_ ), .Z(_101_ ) );
BUF_X1 _542_ ( .A(_064_ ), .Z(_009_ ) );
BUF_X1 _543_ ( .A(\count[2] ), .Z(_128_ ) );
BUF_X1 _544_ ( .A(_047_ ), .Z(_102_ ) );
BUF_X1 _545_ ( .A(_065_ ), .Z(_010_ ) );
BUF_X1 _546_ ( .A(_048_ ), .Z(_103_ ) );
BUF_X1 _547_ ( .A(_066_ ), .Z(_011_ ) );
BUF_X1 _548_ ( .A(\count[3] ), .Z(_129_ ) );
BUF_X1 _549_ ( .A(\count[4] ), .Z(_130_ ) );
BUF_X1 _550_ ( .A(_049_ ), .Z(_104_ ) );
BUF_X1 _551_ ( .A(_067_ ), .Z(_012_ ) );
BUF_X1 _552_ ( .A(_050_ ), .Z(_105_ ) );
BUF_X1 _553_ ( .A(_068_ ), .Z(_013_ ) );
BUF_X1 _554_ ( .A(\count[5] ), .Z(_131_ ) );
BUF_X1 _555_ ( .A(\count[6] ), .Z(_132_ ) );
BUF_X1 _556_ ( .A(_051_ ), .Z(_106_ ) );
BUF_X1 _557_ ( .A(_069_ ), .Z(_014_ ) );
BUF_X1 _558_ ( .A(_052_ ), .Z(_107_ ) );
BUF_X1 _559_ ( .A(_070_ ), .Z(_015_ ) );
DFF_X1 _560_ ( .CK(clk ), .D(_033_ ), .Q(\state[0] ), .QN(_036_ ) );
DFF_X1 _561_ ( .CK(clk ), .D(_034_ ), .Q(\state[1] ), .QN(_054_ ) );
DFF_X1 _562_ ( .CK(clk ), .D(_035_ ), .Q(\state[2] ), .QN(_053_ ) );
DFF_X1 _563_ ( .CK(clk ), .D(_008_ ), .Q(\count[0] ), .QN(_045_ ) );
DFF_X1 _564_ ( .CK(clk ), .D(_009_ ), .Q(\count[1] ), .QN(_046_ ) );
DFF_X1 _565_ ( .CK(clk ), .D(_010_ ), .Q(\count[2] ), .QN(_047_ ) );
DFF_X1 _566_ ( .CK(clk ), .D(_011_ ), .Q(\count[3] ), .QN(_048_ ) );
DFF_X1 _567_ ( .CK(clk ), .D(_012_ ), .Q(\count[4] ), .QN(_049_ ) );
DFF_X1 _568_ ( .CK(clk ), .D(_013_ ), .Q(\count[5] ), .QN(_050_ ) );
DFF_X1 _569_ ( .CK(clk ), .D(_014_ ), .Q(\count[6] ), .QN(_051_ ) );
DFF_X1 _570_ ( .CK(clk ), .D(_015_ ), .Q(\count[7] ), .QN(_052_ ) );
DFF_X1 _571_ ( .CK(clk ), .D(_000_ ), .Q(\buff[0] ), .QN(_037_ ) );
DFF_X1 _572_ ( .CK(clk ), .D(_001_ ), .Q(\buff[1] ), .QN(_038_ ) );
DFF_X1 _573_ ( .CK(clk ), .D(_002_ ), .Q(\buff[2] ), .QN(_039_ ) );
DFF_X1 _574_ ( .CK(clk ), .D(_003_ ), .Q(\buff[3] ), .QN(_040_ ) );
DFF_X1 _575_ ( .CK(clk ), .D(_004_ ), .Q(\buff[4] ), .QN(_041_ ) );
DFF_X1 _576_ ( .CK(clk ), .D(_005_ ), .Q(\buff[5] ), .QN(_042_ ) );
DFF_X1 _577_ ( .CK(clk ), .D(_006_ ), .Q(\buff[6] ), .QN(_043_ ) );
DFF_X1 _578_ ( .CK(clk ), .D(_007_ ), .Q(\buff[7] ), .QN(_044_ ) );
DFF_X1 _579_ ( .CK(clk ), .D(_017_ ), .Q(\ps2_value[0] ), .QN(_281_ ) );
DFF_X1 _580_ ( .CK(clk ), .D(_024_ ), .Q(\ps2_value[1] ), .QN(_282_ ) );
DFF_X1 _581_ ( .CK(clk ), .D(_025_ ), .Q(\ps2_value[2] ), .QN(_283_ ) );
DFF_X1 _582_ ( .CK(clk ), .D(_026_ ), .Q(\ps2_value[3] ), .QN(_284_ ) );
DFF_X1 _583_ ( .CK(clk ), .D(_027_ ), .Q(\ps2_value[4] ), .QN(_285_ ) );
DFF_X1 _584_ ( .CK(clk ), .D(_028_ ), .Q(\ps2_value[5] ), .QN(_286_ ) );
DFF_X1 _585_ ( .CK(clk ), .D(_029_ ), .Q(\ps2_value[6] ), .QN(_287_ ) );
DFF_X1 _586_ ( .CK(clk ), .D(_030_ ), .Q(\ps2_value[7] ), .QN(_288_ ) );
DFF_X1 _587_ ( .CK(clk ), .D(_031_ ), .Q(\ps2_value[8] ), .QN(_289_ ) );
DFF_X1 _588_ ( .CK(clk ), .D(_032_ ), .Q(\ps2_value[9] ), .QN(_290_ ) );
DFF_X1 _589_ ( .CK(clk ), .D(_018_ ), .Q(\ps2_value[10] ), .QN(_291_ ) );
DFF_X1 _590_ ( .CK(clk ), .D(_019_ ), .Q(\ps2_value[11] ), .QN(_292_ ) );
DFF_X1 _591_ ( .CK(clk ), .D(_020_ ), .Q(\ps2_value[12] ), .QN(_293_ ) );
DFF_X1 _592_ ( .CK(clk ), .D(_021_ ), .Q(\ps2_value[13] ), .QN(_294_ ) );
DFF_X1 _593_ ( .CK(clk ), .D(_022_ ), .Q(\ps2_value[14] ), .QN(_295_ ) );
DFF_X1 _594_ ( .CK(clk ), .D(_023_ ), .Q(\ps2_value[15] ), .QN(_296_ ) );
DFF_X1 _595_ ( .CK(clk ), .D(_016_ ), .Q(flag_temp ), .QN(_297_ ) );
LOGIC0_X1 \ScanCodeToASCII_init/_1_ ( .Z(\ScanCodeToASCII_init/_0_ ) );
BUF_X1 \ScanCodeToASCII_init/_2_ ( .A(\ScanCodeToASCII_init/_0_ ), .Z(\ascii_code[0] ) );
BUF_X1 \ScanCodeToASCII_init/_3_ ( .A(\ScanCodeToASCII_init/_0_ ), .Z(\ascii_code[1] ) );
BUF_X1 \ScanCodeToASCII_init/_4_ ( .A(\ScanCodeToASCII_init/_0_ ), .Z(\ascii_code[2] ) );
BUF_X1 \ScanCodeToASCII_init/_5_ ( .A(\ScanCodeToASCII_init/_0_ ), .Z(\ascii_code[3] ) );
BUF_X1 \ScanCodeToASCII_init/_6_ ( .A(\ScanCodeToASCII_init/_0_ ), .Z(\ascii_code[4] ) );
BUF_X1 \ScanCodeToASCII_init/_7_ ( .A(\ScanCodeToASCII_init/_0_ ), .Z(\ascii_code[5] ) );
BUF_X1 \ScanCodeToASCII_init/_8_ ( .A(\ScanCodeToASCII_init/_0_ ), .Z(\ascii_code[6] ) );
BUF_X1 \ScanCodeToASCII_init/_9_ ( .A(\ScanCodeToASCII_init/_0_ ), .Z(\ascii_code[7] ) );
INV_X1 \ps2_keyboard_init/_172_ ( .A(\ps2_keyboard_init/_162_ ), .ZN(\ps2_keyboard_init/_131_ ) );
NOR2_X4 \ps2_keyboard_init/_173_ ( .A1(\ps2_keyboard_init/_131_ ), .A2(\ps2_keyboard_init/_161_ ), .ZN(\ps2_keyboard_init/_132_ ) );
INV_X1 \ps2_keyboard_init/_174_ ( .A(\ps2_keyboard_init/_094_ ), .ZN(\ps2_keyboard_init/_133_ ) );
NOR2_X1 \ps2_keyboard_init/_175_ ( .A1(\ps2_keyboard_init/_133_ ), .A2(\ps2_keyboard_init/_095_ ), .ZN(\ps2_keyboard_init/_134_ ) );
NAND2_X1 \ps2_keyboard_init/_176_ ( .A1(\ps2_keyboard_init/_132_ ), .A2(\ps2_keyboard_init/_134_ ), .ZN(\ps2_keyboard_init/_135_ ) );
INV_X1 \ps2_keyboard_init/_177_ ( .A(\ps2_keyboard_init/_096_ ), .ZN(\ps2_keyboard_init/_136_ ) );
INV_X1 \ps2_keyboard_init/_178_ ( .A(\ps2_keyboard_init/_164_ ), .ZN(\ps2_keyboard_init/_137_ ) );
NAND3_X1 \ps2_keyboard_init/_179_ ( .A1(\ps2_keyboard_init/_136_ ), .A2(\ps2_keyboard_init/_137_ ), .A3(\ps2_keyboard_init/_097_ ), .ZN(\ps2_keyboard_init/_138_ ) );
NOR2_X1 \ps2_keyboard_init/_180_ ( .A1(\ps2_keyboard_init/_135_ ), .A2(\ps2_keyboard_init/_138_ ), .ZN(\ps2_keyboard_init/_139_ ) );
MUX2_X1 \ps2_keyboard_init/_181_ ( .A(\ps2_keyboard_init/_093_ ), .B(\ps2_keyboard_init/_163_ ), .S(\ps2_keyboard_init/_139_ ), .Z(\ps2_keyboard_init/_051_ ) );
NOR3_X1 \ps2_keyboard_init/_182_ ( .A1(\ps2_keyboard_init/_094_ ), .A2(\ps2_keyboard_init/_095_ ), .A3(\ps2_keyboard_init/_164_ ), .ZN(\ps2_keyboard_init/_140_ ) );
INV_X1 \ps2_keyboard_init/_183_ ( .A(\ps2_keyboard_init/_097_ ), .ZN(\ps2_keyboard_init/_141_ ) );
NOR2_X1 \ps2_keyboard_init/_184_ ( .A1(\ps2_keyboard_init/_141_ ), .A2(\ps2_keyboard_init/_096_ ), .ZN(\ps2_keyboard_init/_142_ ) );
NAND3_X1 \ps2_keyboard_init/_185_ ( .A1(\ps2_keyboard_init/_140_ ), .A2(\ps2_keyboard_init/_132_ ), .A3(\ps2_keyboard_init/_142_ ), .ZN(\ps2_keyboard_init/_143_ ) );
MUX2_X1 \ps2_keyboard_init/_186_ ( .A(\ps2_keyboard_init/_163_ ), .B(\ps2_keyboard_init/_092_ ), .S(\ps2_keyboard_init/_143_ ), .Z(\ps2_keyboard_init/_050_ ) );
NOR3_X1 \ps2_keyboard_init/_187_ ( .A1(\ps2_keyboard_init/_136_ ), .A2(\ps2_keyboard_init/_097_ ), .A3(\ps2_keyboard_init/_164_ ), .ZN(\ps2_keyboard_init/_144_ ) );
INV_X1 \ps2_keyboard_init/_188_ ( .A(\ps2_keyboard_init/_144_ ), .ZN(\ps2_keyboard_init/_145_ ) );
AND2_X1 \ps2_keyboard_init/_189_ ( .A1(\ps2_keyboard_init/_094_ ), .A2(\ps2_keyboard_init/_095_ ), .ZN(\ps2_keyboard_init/_146_ ) );
NAND2_X1 \ps2_keyboard_init/_190_ ( .A1(\ps2_keyboard_init/_132_ ), .A2(\ps2_keyboard_init/_146_ ), .ZN(\ps2_keyboard_init/_147_ ) );
NOR2_X1 \ps2_keyboard_init/_191_ ( .A1(\ps2_keyboard_init/_145_ ), .A2(\ps2_keyboard_init/_147_ ), .ZN(\ps2_keyboard_init/_148_ ) );
MUX2_X1 \ps2_keyboard_init/_192_ ( .A(\ps2_keyboard_init/_091_ ), .B(\ps2_keyboard_init/_163_ ), .S(\ps2_keyboard_init/_148_ ), .Z(\ps2_keyboard_init/_049_ ) );
AND3_X1 \ps2_keyboard_init/_193_ ( .A1(\ps2_keyboard_init/_132_ ), .A2(\ps2_keyboard_init/_096_ ), .A3(\ps2_keyboard_init/_141_ ), .ZN(\ps2_keyboard_init/_149_ ) );
AND3_X1 \ps2_keyboard_init/_194_ ( .A1(\ps2_keyboard_init/_133_ ), .A2(\ps2_keyboard_init/_137_ ), .A3(\ps2_keyboard_init/_095_ ), .ZN(\ps2_keyboard_init/_150_ ) );
NAND2_X1 \ps2_keyboard_init/_195_ ( .A1(\ps2_keyboard_init/_149_ ), .A2(\ps2_keyboard_init/_150_ ), .ZN(\ps2_keyboard_init/_151_ ) );
MUX2_X1 \ps2_keyboard_init/_196_ ( .A(\ps2_keyboard_init/_163_ ), .B(\ps2_keyboard_init/_090_ ), .S(\ps2_keyboard_init/_151_ ), .Z(\ps2_keyboard_init/_048_ ) );
NOR2_X1 \ps2_keyboard_init/_197_ ( .A1(\ps2_keyboard_init/_145_ ), .A2(\ps2_keyboard_init/_135_ ), .ZN(\ps2_keyboard_init/_152_ ) );
MUX2_X1 \ps2_keyboard_init/_198_ ( .A(\ps2_keyboard_init/_089_ ), .B(\ps2_keyboard_init/_163_ ), .S(\ps2_keyboard_init/_152_ ), .Z(\ps2_keyboard_init/_047_ ) );
NAND2_X1 \ps2_keyboard_init/_199_ ( .A1(\ps2_keyboard_init/_149_ ), .A2(\ps2_keyboard_init/_140_ ), .ZN(\ps2_keyboard_init/_153_ ) );
MUX2_X1 \ps2_keyboard_init/_200_ ( .A(\ps2_keyboard_init/_163_ ), .B(\ps2_keyboard_init/_088_ ), .S(\ps2_keyboard_init/_153_ ), .Z(\ps2_keyboard_init/_046_ ) );
NOR2_X1 \ps2_keyboard_init/_201_ ( .A1(\ps2_keyboard_init/_096_ ), .A2(\ps2_keyboard_init/_097_ ), .ZN(\ps2_keyboard_init/_154_ ) );
AND2_X1 \ps2_keyboard_init/_202_ ( .A1(\ps2_keyboard_init/_132_ ), .A2(\ps2_keyboard_init/_154_ ), .ZN(\ps2_keyboard_init/_155_ ) );
AND3_X1 \ps2_keyboard_init/_203_ ( .A1(\ps2_keyboard_init/_137_ ), .A2(\ps2_keyboard_init/_094_ ), .A3(\ps2_keyboard_init/_095_ ), .ZN(\ps2_keyboard_init/_156_ ) );
NAND2_X1 \ps2_keyboard_init/_204_ ( .A1(\ps2_keyboard_init/_155_ ), .A2(\ps2_keyboard_init/_156_ ), .ZN(\ps2_keyboard_init/_157_ ) );
MUX2_X1 \ps2_keyboard_init/_205_ ( .A(\ps2_keyboard_init/_163_ ), .B(\ps2_keyboard_init/_087_ ), .S(\ps2_keyboard_init/_157_ ), .Z(\ps2_keyboard_init/_045_ ) );
NAND2_X1 \ps2_keyboard_init/_206_ ( .A1(\ps2_keyboard_init/_155_ ), .A2(\ps2_keyboard_init/_150_ ), .ZN(\ps2_keyboard_init/_158_ ) );
MUX2_X1 \ps2_keyboard_init/_207_ ( .A(\ps2_keyboard_init/_163_ ), .B(\ps2_keyboard_init/_086_ ), .S(\ps2_keyboard_init/_158_ ), .Z(\ps2_keyboard_init/_044_ ) );
NOR3_X1 \ps2_keyboard_init/_208_ ( .A1(\ps2_keyboard_init/_133_ ), .A2(\ps2_keyboard_init/_095_ ), .A3(\ps2_keyboard_init/_164_ ), .ZN(\ps2_keyboard_init/_159_ ) );
NAND2_X1 \ps2_keyboard_init/_209_ ( .A1(\ps2_keyboard_init/_155_ ), .A2(\ps2_keyboard_init/_159_ ), .ZN(\ps2_keyboard_init/_160_ ) );
MUX2_X1 \ps2_keyboard_init/_210_ ( .A(\ps2_keyboard_init/_163_ ), .B(\ps2_keyboard_init/_085_ ), .S(\ps2_keyboard_init/_160_ ), .Z(\ps2_keyboard_init/_043_ ) );
NAND2_X1 \ps2_keyboard_init/_211_ ( .A1(\ps2_keyboard_init/_155_ ), .A2(\ps2_keyboard_init/_140_ ), .ZN(\ps2_keyboard_init/_098_ ) );
MUX2_X1 \ps2_keyboard_init/_212_ ( .A(\ps2_keyboard_init/_163_ ), .B(\ps2_keyboard_init/_084_ ), .S(\ps2_keyboard_init/_098_ ), .Z(\ps2_keyboard_init/_042_ ) );
XNOR2_X2 \ps2_keyboard_init/_213_ ( .A(\ps2_keyboard_init/_092_ ), .B(\ps2_keyboard_init/_091_ ), .ZN(\ps2_keyboard_init/_099_ ) );
XNOR2_X2 \ps2_keyboard_init/_214_ ( .A(\ps2_keyboard_init/_090_ ), .B(\ps2_keyboard_init/_089_ ), .ZN(\ps2_keyboard_init/_100_ ) );
XOR2_X1 \ps2_keyboard_init/_215_ ( .A(\ps2_keyboard_init/_099_ ), .B(\ps2_keyboard_init/_100_ ), .Z(\ps2_keyboard_init/_101_ ) );
XOR2_X2 \ps2_keyboard_init/_216_ ( .A(\ps2_keyboard_init/_086_ ), .B(\ps2_keyboard_init/_085_ ), .Z(\ps2_keyboard_init/_102_ ) );
XNOR2_X2 \ps2_keyboard_init/_217_ ( .A(\ps2_keyboard_init/_088_ ), .B(\ps2_keyboard_init/_087_ ), .ZN(\ps2_keyboard_init/_103_ ) );
XNOR2_X2 \ps2_keyboard_init/_218_ ( .A(\ps2_keyboard_init/_102_ ), .B(\ps2_keyboard_init/_103_ ), .ZN(\ps2_keyboard_init/_104_ ) );
XNOR2_X2 \ps2_keyboard_init/_219_ ( .A(\ps2_keyboard_init/_101_ ), .B(\ps2_keyboard_init/_104_ ), .ZN(\ps2_keyboard_init/_105_ ) );
XNOR2_X2 \ps2_keyboard_init/_220_ ( .A(\ps2_keyboard_init/_105_ ), .B(\ps2_keyboard_init/_093_ ), .ZN(\ps2_keyboard_init/_106_ ) );
AND2_X1 \ps2_keyboard_init/_221_ ( .A1(\ps2_keyboard_init/_132_ ), .A2(\ps2_keyboard_init/_142_ ), .ZN(\ps2_keyboard_init/_107_ ) );
AND2_X1 \ps2_keyboard_init/_222_ ( .A1(\ps2_keyboard_init/_133_ ), .A2(\ps2_keyboard_init/_095_ ), .ZN(\ps2_keyboard_init/_108_ ) );
AND2_X1 \ps2_keyboard_init/_223_ ( .A1(\ps2_keyboard_init/_107_ ), .A2(\ps2_keyboard_init/_108_ ), .ZN(\ps2_keyboard_init/_109_ ) );
INV_X1 \ps2_keyboard_init/_224_ ( .A(\ps2_keyboard_init/_109_ ), .ZN(\ps2_keyboard_init/_110_ ) );
NOR2_X1 \ps2_keyboard_init/_225_ ( .A1(\ps2_keyboard_init/_110_ ), .A2(\ps2_keyboard_init/_084_ ), .ZN(\ps2_keyboard_init/_111_ ) );
AND2_X2 \ps2_keyboard_init/_226_ ( .A1(\ps2_keyboard_init/_111_ ), .A2(\ps2_keyboard_init/_163_ ), .ZN(\ps2_keyboard_init/_112_ ) );
AND3_X1 \ps2_keyboard_init/_227_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_066_ ), .A3(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_113_ ) );
NAND2_X4 \ps2_keyboard_init/_228_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_114_ ) );
AOI211_X2 \ps2_keyboard_init/_229_ ( .A(\ps2_keyboard_init/_164_ ), .B(\ps2_keyboard_init/_113_ ), .C1(\ps2_keyboard_init/_065_ ), .C2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_056_ ) );
AND3_X1 \ps2_keyboard_init/_230_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_068_ ), .A3(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_115_ ) );
AOI211_X2 \ps2_keyboard_init/_231_ ( .A(\ps2_keyboard_init/_164_ ), .B(\ps2_keyboard_init/_115_ ), .C1(\ps2_keyboard_init/_067_ ), .C2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_057_ ) );
AND3_X1 \ps2_keyboard_init/_232_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_070_ ), .A3(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_116_ ) );
AOI211_X2 \ps2_keyboard_init/_233_ ( .A(\ps2_keyboard_init/_164_ ), .B(\ps2_keyboard_init/_116_ ), .C1(\ps2_keyboard_init/_069_ ), .C2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_058_ ) );
AND3_X1 \ps2_keyboard_init/_234_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_072_ ), .A3(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_117_ ) );
AOI211_X2 \ps2_keyboard_init/_235_ ( .A(\ps2_keyboard_init/_164_ ), .B(\ps2_keyboard_init/_117_ ), .C1(\ps2_keyboard_init/_071_ ), .C2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_059_ ) );
AND3_X1 \ps2_keyboard_init/_236_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_074_ ), .A3(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_118_ ) );
AOI211_X2 \ps2_keyboard_init/_237_ ( .A(\ps2_keyboard_init/_164_ ), .B(\ps2_keyboard_init/_118_ ), .C1(\ps2_keyboard_init/_073_ ), .C2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_060_ ) );
AND3_X1 \ps2_keyboard_init/_238_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_076_ ), .A3(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_119_ ) );
AOI211_X2 \ps2_keyboard_init/_239_ ( .A(\ps2_keyboard_init/_164_ ), .B(\ps2_keyboard_init/_119_ ), .C1(\ps2_keyboard_init/_075_ ), .C2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_061_ ) );
AND3_X1 \ps2_keyboard_init/_240_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_078_ ), .A3(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_120_ ) );
AOI211_X2 \ps2_keyboard_init/_241_ ( .A(\ps2_keyboard_init/_164_ ), .B(\ps2_keyboard_init/_120_ ), .C1(\ps2_keyboard_init/_077_ ), .C2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_062_ ) );
AND3_X1 \ps2_keyboard_init/_242_ ( .A1(\ps2_keyboard_init/_106_ ), .A2(\ps2_keyboard_init/_080_ ), .A3(\ps2_keyboard_init/_112_ ), .ZN(\ps2_keyboard_init/_121_ ) );
AOI211_X2 \ps2_keyboard_init/_243_ ( .A(\ps2_keyboard_init/_164_ ), .B(\ps2_keyboard_init/_121_ ), .C1(\ps2_keyboard_init/_079_ ), .C2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_063_ ) );
AOI21_X1 \ps2_keyboard_init/_244_ ( .A(\ps2_keyboard_init/_109_ ), .B1(\ps2_keyboard_init/_094_ ), .B2(\ps2_keyboard_init/_132_ ), .ZN(\ps2_keyboard_init/_122_ ) );
OAI21_X1 \ps2_keyboard_init/_245_ ( .A(\ps2_keyboard_init/_081_ ), .B1(\ps2_keyboard_init/_131_ ), .B2(\ps2_keyboard_init/_161_ ), .ZN(\ps2_keyboard_init/_123_ ) );
AND3_X1 \ps2_keyboard_init/_246_ ( .A1(\ps2_keyboard_init/_122_ ), .A2(\ps2_keyboard_init/_137_ ), .A3(\ps2_keyboard_init/_123_ ), .ZN(\ps2_keyboard_init/_052_ ) );
NAND2_X1 \ps2_keyboard_init/_247_ ( .A1(\ps2_keyboard_init/_122_ ), .A2(\ps2_keyboard_init/_095_ ), .ZN(\ps2_keyboard_init/_124_ ) );
AOI21_X1 \ps2_keyboard_init/_248_ ( .A(\ps2_keyboard_init/_164_ ), .B1(\ps2_keyboard_init/_124_ ), .B2(\ps2_keyboard_init/_135_ ), .ZN(\ps2_keyboard_init/_053_ ) );
AND3_X1 \ps2_keyboard_init/_249_ ( .A1(\ps2_keyboard_init/_132_ ), .A2(\ps2_keyboard_init/_096_ ), .A3(\ps2_keyboard_init/_146_ ), .ZN(\ps2_keyboard_init/_125_ ) );
INV_X1 \ps2_keyboard_init/_250_ ( .A(\ps2_keyboard_init/_125_ ), .ZN(\ps2_keyboard_init/_126_ ) );
AOI21_X1 \ps2_keyboard_init/_251_ ( .A(\ps2_keyboard_init/_164_ ), .B1(\ps2_keyboard_init/_147_ ), .B2(\ps2_keyboard_init/_136_ ), .ZN(\ps2_keyboard_init/_127_ ) );
AND2_X1 \ps2_keyboard_init/_252_ ( .A1(\ps2_keyboard_init/_126_ ), .A2(\ps2_keyboard_init/_127_ ), .ZN(\ps2_keyboard_init/_054_ ) );
AOI221_X4 \ps2_keyboard_init/_253_ ( .A(\ps2_keyboard_init/_164_ ), .B1(\ps2_keyboard_init/_107_ ), .B2(\ps2_keyboard_init/_108_ ), .C1(\ps2_keyboard_init/_126_ ), .C2(\ps2_keyboard_init/_082_ ), .ZN(\ps2_keyboard_init/_128_ ) );
OR3_X1 \ps2_keyboard_init/_254_ ( .A1(\ps2_keyboard_init/_147_ ), .A2(\ps2_keyboard_init/_136_ ), .A3(\ps2_keyboard_init/_082_ ), .ZN(\ps2_keyboard_init/_129_ ) );
AND2_X1 \ps2_keyboard_init/_255_ ( .A1(\ps2_keyboard_init/_128_ ), .A2(\ps2_keyboard_init/_129_ ), .ZN(\ps2_keyboard_init/_055_ ) );
OAI21_X2 \ps2_keyboard_init/_256_ ( .A(\ps2_keyboard_init/_137_ ), .B1(\ps2_keyboard_init/_114_ ), .B2(\ps2_keyboard_init/_083_ ), .ZN(\ps2_keyboard_init/_130_ ) );
AOI21_X1 \ps2_keyboard_init/_257_ ( .A(\ps2_keyboard_init/_130_ ), .B1(\ps2_keyboard_init/_083_ ), .B2(\ps2_keyboard_init/_114_ ), .ZN(\ps2_keyboard_init/_064_ ) );
BUF_X1 \ps2_keyboard_init/_258_ ( .A(\ps2_keyboard_init/ps2_clk_sync[1] ), .Z(\ps2_keyboard_init/_161_ ) );
BUF_X1 \ps2_keyboard_init/_259_ ( .A(\ps2_keyboard_init/ps2_clk_sync[2] ), .Z(\ps2_keyboard_init/_162_ ) );
BUF_X1 \ps2_keyboard_init/_260_ ( .A(\ps2_keyboard_init/count[2] ), .Z(\ps2_keyboard_init/_096_ ) );
BUF_X1 \ps2_keyboard_init/_261_ ( .A(\ps2_keyboard_init/count[3] ), .Z(\ps2_keyboard_init/_097_ ) );
BUF_X1 \ps2_keyboard_init/_262_ ( .A(\ps2_keyboard_init/count[0] ), .Z(\ps2_keyboard_init/_094_ ) );
BUF_X1 \ps2_keyboard_init/_263_ ( .A(\ps2_keyboard_init/count[1] ), .Z(\ps2_keyboard_init/_095_ ) );
BUF_X1 \ps2_keyboard_init/_264_ ( .A(ps2_data ), .Z(\ps2_keyboard_init/_163_ ) );
BUF_X1 \ps2_keyboard_init/_265_ ( .A(\ps2_keyboard_init/buffer[9] ), .Z(\ps2_keyboard_init/_093_ ) );
BUF_X1 \ps2_keyboard_init/_266_ ( .A(rst_n ), .Z(\ps2_keyboard_init/_164_ ) );
BUF_X1 \ps2_keyboard_init/_267_ ( .A(\ps2_keyboard_init/_051_ ), .Z(\ps2_keyboard_init/_009_ ) );
BUF_X1 \ps2_keyboard_init/_268_ ( .A(\ps2_keyboard_init/buffer[8] ), .Z(\ps2_keyboard_init/_092_ ) );
BUF_X1 \ps2_keyboard_init/_269_ ( .A(\ps2_keyboard_init/_050_ ), .Z(\ps2_keyboard_init/_008_ ) );
BUF_X1 \ps2_keyboard_init/_270_ ( .A(\ps2_keyboard_init/buffer[7] ), .Z(\ps2_keyboard_init/_091_ ) );
BUF_X1 \ps2_keyboard_init/_271_ ( .A(\ps2_keyboard_init/_049_ ), .Z(\ps2_keyboard_init/_007_ ) );
BUF_X1 \ps2_keyboard_init/_272_ ( .A(\ps2_keyboard_init/buffer[6] ), .Z(\ps2_keyboard_init/_090_ ) );
BUF_X1 \ps2_keyboard_init/_273_ ( .A(\ps2_keyboard_init/_048_ ), .Z(\ps2_keyboard_init/_006_ ) );
BUF_X1 \ps2_keyboard_init/_274_ ( .A(\ps2_keyboard_init/buffer[5] ), .Z(\ps2_keyboard_init/_089_ ) );
BUF_X1 \ps2_keyboard_init/_275_ ( .A(\ps2_keyboard_init/_047_ ), .Z(\ps2_keyboard_init/_005_ ) );
BUF_X1 \ps2_keyboard_init/_276_ ( .A(\ps2_keyboard_init/buffer[4] ), .Z(\ps2_keyboard_init/_088_ ) );
BUF_X1 \ps2_keyboard_init/_277_ ( .A(\ps2_keyboard_init/_046_ ), .Z(\ps2_keyboard_init/_004_ ) );
BUF_X1 \ps2_keyboard_init/_278_ ( .A(\ps2_keyboard_init/buffer[3] ), .Z(\ps2_keyboard_init/_087_ ) );
BUF_X1 \ps2_keyboard_init/_279_ ( .A(\ps2_keyboard_init/_045_ ), .Z(\ps2_keyboard_init/_003_ ) );
BUF_X1 \ps2_keyboard_init/_280_ ( .A(\ps2_keyboard_init/buffer[2] ), .Z(\ps2_keyboard_init/_086_ ) );
BUF_X1 \ps2_keyboard_init/_281_ ( .A(\ps2_keyboard_init/_044_ ), .Z(\ps2_keyboard_init/_002_ ) );
BUF_X1 \ps2_keyboard_init/_282_ ( .A(\ps2_keyboard_init/buffer[1] ), .Z(\ps2_keyboard_init/_085_ ) );
BUF_X1 \ps2_keyboard_init/_283_ ( .A(\ps2_keyboard_init/_043_ ), .Z(\ps2_keyboard_init/_001_ ) );
BUF_X1 \ps2_keyboard_init/_284_ ( .A(\ps2_keyboard_init/buffer[0] ), .Z(\ps2_keyboard_init/_084_ ) );
BUF_X1 \ps2_keyboard_init/_285_ ( .A(\ps2_keyboard_init/_042_ ), .Z(\ps2_keyboard_init/_000_ ) );
BUF_X1 \ps2_keyboard_init/_286_ ( .A(\ps2_keyboard_init/_023_ ), .Z(\ps2_keyboard_init/_065_ ) );
BUF_X1 \ps2_keyboard_init/_287_ ( .A(\ps2_keyboard_init/_024_ ), .Z(\ps2_keyboard_init/_066_ ) );
BUF_X1 \ps2_keyboard_init/_288_ ( .A(\ps2_keyboard_init/_056_ ), .Z(\ps2_keyboard_init/_014_ ) );
BUF_X1 \ps2_keyboard_init/_289_ ( .A(\ps2_keyboard_init/_025_ ), .Z(\ps2_keyboard_init/_067_ ) );
BUF_X1 \ps2_keyboard_init/_290_ ( .A(\ps2_keyboard_init/_026_ ), .Z(\ps2_keyboard_init/_068_ ) );
BUF_X1 \ps2_keyboard_init/_291_ ( .A(\ps2_keyboard_init/_057_ ), .Z(\ps2_keyboard_init/_015_ ) );
BUF_X1 \ps2_keyboard_init/_292_ ( .A(\ps2_keyboard_init/_027_ ), .Z(\ps2_keyboard_init/_069_ ) );
BUF_X1 \ps2_keyboard_init/_293_ ( .A(\ps2_keyboard_init/_028_ ), .Z(\ps2_keyboard_init/_070_ ) );
BUF_X1 \ps2_keyboard_init/_294_ ( .A(\ps2_keyboard_init/_058_ ), .Z(\ps2_keyboard_init/_016_ ) );
BUF_X1 \ps2_keyboard_init/_295_ ( .A(\ps2_keyboard_init/_029_ ), .Z(\ps2_keyboard_init/_071_ ) );
BUF_X1 \ps2_keyboard_init/_296_ ( .A(\ps2_keyboard_init/_030_ ), .Z(\ps2_keyboard_init/_072_ ) );
BUF_X1 \ps2_keyboard_init/_297_ ( .A(\ps2_keyboard_init/_059_ ), .Z(\ps2_keyboard_init/_017_ ) );
BUF_X1 \ps2_keyboard_init/_298_ ( .A(\ps2_keyboard_init/_031_ ), .Z(\ps2_keyboard_init/_073_ ) );
BUF_X1 \ps2_keyboard_init/_299_ ( .A(\ps2_keyboard_init/_032_ ), .Z(\ps2_keyboard_init/_074_ ) );
BUF_X1 \ps2_keyboard_init/_300_ ( .A(\ps2_keyboard_init/_060_ ), .Z(\ps2_keyboard_init/_018_ ) );
BUF_X1 \ps2_keyboard_init/_301_ ( .A(\ps2_keyboard_init/_033_ ), .Z(\ps2_keyboard_init/_075_ ) );
BUF_X1 \ps2_keyboard_init/_302_ ( .A(\ps2_keyboard_init/_034_ ), .Z(\ps2_keyboard_init/_076_ ) );
BUF_X1 \ps2_keyboard_init/_303_ ( .A(\ps2_keyboard_init/_061_ ), .Z(\ps2_keyboard_init/_019_ ) );
BUF_X1 \ps2_keyboard_init/_304_ ( .A(\ps2_keyboard_init/_035_ ), .Z(\ps2_keyboard_init/_077_ ) );
BUF_X1 \ps2_keyboard_init/_305_ ( .A(\ps2_keyboard_init/_036_ ), .Z(\ps2_keyboard_init/_078_ ) );
BUF_X1 \ps2_keyboard_init/_306_ ( .A(\ps2_keyboard_init/_062_ ), .Z(\ps2_keyboard_init/_020_ ) );
BUF_X1 \ps2_keyboard_init/_307_ ( .A(\ps2_keyboard_init/_037_ ), .Z(\ps2_keyboard_init/_079_ ) );
BUF_X1 \ps2_keyboard_init/_308_ ( .A(\ps2_keyboard_init/_038_ ), .Z(\ps2_keyboard_init/_080_ ) );
BUF_X1 \ps2_keyboard_init/_309_ ( .A(\ps2_keyboard_init/_063_ ), .Z(\ps2_keyboard_init/_021_ ) );
BUF_X1 \ps2_keyboard_init/_310_ ( .A(\ps2_keyboard_init/_039_ ), .Z(\ps2_keyboard_init/_081_ ) );
BUF_X1 \ps2_keyboard_init/_311_ ( .A(\ps2_keyboard_init/_052_ ), .Z(\ps2_keyboard_init/_010_ ) );
BUF_X1 \ps2_keyboard_init/_312_ ( .A(\ps2_keyboard_init/_053_ ), .Z(\ps2_keyboard_init/_011_ ) );
BUF_X1 \ps2_keyboard_init/_313_ ( .A(\ps2_keyboard_init/_054_ ), .Z(\ps2_keyboard_init/_012_ ) );
BUF_X1 \ps2_keyboard_init/_314_ ( .A(\ps2_keyboard_init/_040_ ), .Z(\ps2_keyboard_init/_082_ ) );
BUF_X1 \ps2_keyboard_init/_315_ ( .A(\ps2_keyboard_init/_055_ ), .Z(\ps2_keyboard_init/_013_ ) );
BUF_X1 \ps2_keyboard_init/_316_ ( .A(\ps2_keyboard_init/_041_ ), .Z(\ps2_keyboard_init/_083_ ) );
BUF_X1 \ps2_keyboard_init/_317_ ( .A(\ps2_keyboard_init/_064_ ), .Z(\ps2_keyboard_init/_022_ ) );
DFF_X1 \ps2_keyboard_init/_318_ ( .CK(clk ), .D(\ps2_keyboard_init/_000_ ), .Q(\ps2_keyboard_init/buffer[0] ), .QN(\ps2_keyboard_init/_165_ ) );
DFF_X1 \ps2_keyboard_init/_319_ ( .CK(clk ), .D(\ps2_keyboard_init/_001_ ), .Q(\ps2_keyboard_init/buffer[1] ), .QN(\ps2_keyboard_init/_024_ ) );
DFF_X1 \ps2_keyboard_init/_320_ ( .CK(clk ), .D(\ps2_keyboard_init/_002_ ), .Q(\ps2_keyboard_init/buffer[2] ), .QN(\ps2_keyboard_init/_026_ ) );
DFF_X1 \ps2_keyboard_init/_321_ ( .CK(clk ), .D(\ps2_keyboard_init/_003_ ), .Q(\ps2_keyboard_init/buffer[3] ), .QN(\ps2_keyboard_init/_028_ ) );
DFF_X1 \ps2_keyboard_init/_322_ ( .CK(clk ), .D(\ps2_keyboard_init/_004_ ), .Q(\ps2_keyboard_init/buffer[4] ), .QN(\ps2_keyboard_init/_030_ ) );
DFF_X1 \ps2_keyboard_init/_323_ ( .CK(clk ), .D(\ps2_keyboard_init/_005_ ), .Q(\ps2_keyboard_init/buffer[5] ), .QN(\ps2_keyboard_init/_032_ ) );
DFF_X1 \ps2_keyboard_init/_324_ ( .CK(clk ), .D(\ps2_keyboard_init/_006_ ), .Q(\ps2_keyboard_init/buffer[6] ), .QN(\ps2_keyboard_init/_034_ ) );
DFF_X1 \ps2_keyboard_init/_325_ ( .CK(clk ), .D(\ps2_keyboard_init/_007_ ), .Q(\ps2_keyboard_init/buffer[7] ), .QN(\ps2_keyboard_init/_036_ ) );
DFF_X1 \ps2_keyboard_init/_326_ ( .CK(clk ), .D(\ps2_keyboard_init/_008_ ), .Q(\ps2_keyboard_init/buffer[8] ), .QN(\ps2_keyboard_init/_038_ ) );
DFF_X1 \ps2_keyboard_init/_327_ ( .CK(clk ), .D(\ps2_keyboard_init/_009_ ), .Q(\ps2_keyboard_init/buffer[9] ), .QN(\ps2_keyboard_init/_166_ ) );
DFF_X1 \ps2_keyboard_init/_328_ ( .CK(clk ), .D(\ps2_keyboard_init/_010_ ), .Q(\ps2_keyboard_init/count[0] ), .QN(\ps2_keyboard_init/_039_ ) );
DFF_X1 \ps2_keyboard_init/_329_ ( .CK(clk ), .D(\ps2_keyboard_init/_011_ ), .Q(\ps2_keyboard_init/count[1] ), .QN(\ps2_keyboard_init/_167_ ) );
DFF_X1 \ps2_keyboard_init/_330_ ( .CK(clk ), .D(\ps2_keyboard_init/_012_ ), .Q(\ps2_keyboard_init/count[2] ), .QN(\ps2_keyboard_init/_168_ ) );
DFF_X1 \ps2_keyboard_init/_331_ ( .CK(clk ), .D(\ps2_keyboard_init/_013_ ), .Q(\ps2_keyboard_init/count[3] ), .QN(\ps2_keyboard_init/_040_ ) );
DFF_X1 \ps2_keyboard_init/_332_ ( .CK(clk ), .D(\ps2_keyboard_init/_014_ ), .Q(\data[0] ), .QN(\ps2_keyboard_init/_023_ ) );
DFF_X1 \ps2_keyboard_init/_333_ ( .CK(clk ), .D(\ps2_keyboard_init/_015_ ), .Q(\data[1] ), .QN(\ps2_keyboard_init/_025_ ) );
DFF_X1 \ps2_keyboard_init/_334_ ( .CK(clk ), .D(\ps2_keyboard_init/_016_ ), .Q(\data[2] ), .QN(\ps2_keyboard_init/_027_ ) );
DFF_X1 \ps2_keyboard_init/_335_ ( .CK(clk ), .D(\ps2_keyboard_init/_017_ ), .Q(\data[3] ), .QN(\ps2_keyboard_init/_029_ ) );
DFF_X1 \ps2_keyboard_init/_336_ ( .CK(clk ), .D(\ps2_keyboard_init/_018_ ), .Q(\data[4] ), .QN(\ps2_keyboard_init/_031_ ) );
DFF_X1 \ps2_keyboard_init/_337_ ( .CK(clk ), .D(\ps2_keyboard_init/_019_ ), .Q(\data[5] ), .QN(\ps2_keyboard_init/_033_ ) );
DFF_X1 \ps2_keyboard_init/_338_ ( .CK(clk ), .D(\ps2_keyboard_init/_020_ ), .Q(\data[6] ), .QN(\ps2_keyboard_init/_035_ ) );
DFF_X1 \ps2_keyboard_init/_339_ ( .CK(clk ), .D(\ps2_keyboard_init/_021_ ), .Q(\data[7] ), .QN(\ps2_keyboard_init/_037_ ) );
DFF_X1 \ps2_keyboard_init/_340_ ( .CK(clk ), .D(\ps2_keyboard_init/_022_ ), .Q(flag ), .QN(\ps2_keyboard_init/_041_ ) );
DFF_X1 \ps2_keyboard_init/_341_ ( .CK(clk ), .D(ps2_clk ), .Q(\ps2_keyboard_init/ps2_clk_sync[0] ), .QN(\ps2_keyboard_init/_169_ ) );
DFF_X1 \ps2_keyboard_init/_342_ ( .CK(clk ), .D(\ps2_keyboard_init/ps2_clk_sync[0] ), .Q(\ps2_keyboard_init/ps2_clk_sync[1] ), .QN(\ps2_keyboard_init/_170_ ) );
DFF_X1 \ps2_keyboard_init/_343_ ( .CK(clk ), .D(\ps2_keyboard_init/ps2_clk_sync[1] ), .Q(\ps2_keyboard_init/ps2_clk_sync[2] ), .QN(\ps2_keyboard_init/_171_ ) );
INV_X16 \seg0/_38_ ( .A(\seg0/_00_ ), .ZN(\seg0/_11_ ) );
NOR2_X4 \seg0/_39_ ( .A1(\seg0/_11_ ), .A2(\seg0/_01_ ), .ZN(\seg0/_12_ ) );
AND2_X4 \seg0/_40_ ( .A1(\seg0/_03_ ), .A2(\seg0/_02_ ), .ZN(\seg0/_13_ ) );
AND2_X4 \seg0/_41_ ( .A1(\seg0/_12_ ), .A2(\seg0/_13_ ), .ZN(\seg0/_14_ ) );
NOR2_X4 \seg0/_42_ ( .A1(\seg0/_00_ ), .A2(\seg0/_01_ ), .ZN(\seg0/_15_ ) );
INV_X32 \seg0/_43_ ( .A(\seg0/_02_ ), .ZN(\seg0/_16_ ) );
NOR2_X4 \seg0/_44_ ( .A1(\seg0/_16_ ), .A2(\seg0/_03_ ), .ZN(\seg0/_17_ ) );
AOI21_X4 \seg0/_45_ ( .A(\seg0/_14_ ), .B1(\seg0/_15_ ), .B2(\seg0/_17_ ), .ZN(\seg0/_18_ ) );
AND2_X4 \seg0/_46_ ( .A1(\seg0/_00_ ), .A2(\seg0/_01_ ), .ZN(\seg0/_19_ ) );
AND3_X2 \seg0/_47_ ( .A1(\seg0/_19_ ), .A2(\seg0/_03_ ), .A3(\seg0/_16_ ), .ZN(\seg0/_20_ ) );
NOR2_X4 \seg0/_48_ ( .A1(\seg0/_03_ ), .A2(\seg0/_02_ ), .ZN(\seg0/_21_ ) );
AND2_X1 \seg0/_49_ ( .A1(\seg0/_15_ ), .A2(\seg0/_21_ ), .ZN(\seg0/_22_ ) );
NOR2_X2 \seg0/_50_ ( .A1(\seg0/_20_ ), .A2(\seg0/_22_ ), .ZN(\seg0/_23_ ) );
INV_X1 \seg0/_51_ ( .A(\seg0/_21_ ), .ZN(\seg0/_24_ ) );
INV_X1 \seg0/_52_ ( .A(\seg0/_12_ ), .ZN(\seg0/_25_ ) );
OAI211_X2 \seg0/_53_ ( .A(\seg0/_18_ ), .B(\seg0/_23_ ), .C1(\seg0/_24_ ), .C2(\seg0/_25_ ), .ZN(\seg0/_04_ ) );
INV_X16 \seg0/_54_ ( .A(\seg0/_01_ ), .ZN(\seg0/_26_ ) );
NOR2_X4 \seg0/_55_ ( .A1(\seg0/_26_ ), .A2(\seg0/_00_ ), .ZN(\seg0/_27_ ) );
OAI21_X1 \seg0/_56_ ( .A(\seg0/_17_ ), .B1(\seg0/_12_ ), .B2(\seg0/_27_ ), .ZN(\seg0/_28_ ) );
NAND2_X1 \seg0/_57_ ( .A1(\seg0/_25_ ), .A2(\seg0/_13_ ), .ZN(\seg0/_29_ ) );
NAND3_X1 \seg0/_58_ ( .A1(\seg0/_23_ ), .A2(\seg0/_28_ ), .A3(\seg0/_29_ ), .ZN(\seg0/_05_ ) );
OAI21_X1 \seg0/_59_ ( .A(\seg0/_29_ ), .B1(\seg0/_00_ ), .B2(\seg0/_24_ ), .ZN(\seg0/_06_ ) );
INV_X1 \seg0/_60_ ( .A(\seg0/_17_ ), .ZN(\seg0/_30_ ) );
OR3_X2 \seg0/_61_ ( .A1(\seg0/_30_ ), .A2(\seg0/_12_ ), .A3(\seg0/_27_ ), .ZN(\seg0/_31_ ) );
NAND3_X1 \seg0/_62_ ( .A1(\seg0/_27_ ), .A2(\seg0/_03_ ), .A3(\seg0/_16_ ), .ZN(\seg0/_32_ ) );
NAND2_X1 \seg0/_63_ ( .A1(\seg0/_19_ ), .A2(\seg0/_13_ ), .ZN(\seg0/_33_ ) );
NAND2_X1 \seg0/_64_ ( .A1(\seg0/_21_ ), .A2(\seg0/_26_ ), .ZN(\seg0/_34_ ) );
NAND4_X1 \seg0/_65_ ( .A1(\seg0/_31_ ), .A2(\seg0/_32_ ), .A3(\seg0/_33_ ), .A4(\seg0/_34_ ), .ZN(\seg0/_07_ ) );
OAI22_X1 \seg0/_66_ ( .A1(\seg0/_25_ ), .A2(\seg0/_02_ ), .B1(\seg0/_03_ ), .B2(\seg0/_27_ ), .ZN(\seg0/_08_ ) );
AOI22_X1 \seg0/_67_ ( .A1(\seg0/_12_ ), .A2(\seg0/_13_ ), .B1(\seg0/_15_ ), .B2(\seg0/_21_ ), .ZN(\seg0/_35_ ) );
NAND2_X1 \seg0/_68_ ( .A1(\seg0/_17_ ), .A2(\seg0/_19_ ), .ZN(\seg0/_36_ ) );
OAI211_X2 \seg0/_69_ ( .A(\seg0/_35_ ), .B(\seg0/_36_ ), .C1(\seg0/_15_ ), .C2(\seg0/_24_ ), .ZN(\seg0/_09_ ) );
NAND2_X1 \seg0/_70_ ( .A1(\seg0/_13_ ), .A2(\seg0/_15_ ), .ZN(\seg0/_37_ ) );
NAND3_X1 \seg0/_71_ ( .A1(\seg0/_36_ ), .A2(\seg0/_34_ ), .A3(\seg0/_37_ ), .ZN(\seg0/_10_ ) );
BUF_X1 \seg0/_72_ ( .A(\ps2_value[3] ), .Z(\seg0/_03_ ) );
BUF_X1 \seg0/_73_ ( .A(\ps2_value[2] ), .Z(\seg0/_02_ ) );
BUF_X1 \seg0/_74_ ( .A(\ps2_value[0] ), .Z(\seg0/_00_ ) );
BUF_X1 \seg0/_75_ ( .A(\ps2_value[1] ), .Z(\seg0/_01_ ) );
BUF_X1 \seg0/_76_ ( .A(\seg0/_04_ ), .Z(\value_seg[0] ) );
BUF_X1 \seg0/_77_ ( .A(\seg0/_05_ ), .Z(\value_seg[1] ) );
BUF_X1 \seg0/_78_ ( .A(\seg0/_06_ ), .Z(\value_seg[2] ) );
BUF_X1 \seg0/_79_ ( .A(\seg0/_07_ ), .Z(\value_seg[3] ) );
BUF_X1 \seg0/_80_ ( .A(\seg0/_08_ ), .Z(\value_seg[4] ) );
BUF_X1 \seg0/_81_ ( .A(\seg0/_09_ ), .Z(\value_seg[5] ) );
BUF_X1 \seg0/_82_ ( .A(\seg0/_10_ ), .Z(\value_seg[6] ) );
INV_X16 \seg1/_38_ ( .A(\seg1/_00_ ), .ZN(\seg1/_11_ ) );
NOR2_X4 \seg1/_39_ ( .A1(\seg1/_11_ ), .A2(\seg1/_01_ ), .ZN(\seg1/_12_ ) );
AND2_X4 \seg1/_40_ ( .A1(\seg1/_03_ ), .A2(\seg1/_02_ ), .ZN(\seg1/_13_ ) );
AND2_X4 \seg1/_41_ ( .A1(\seg1/_12_ ), .A2(\seg1/_13_ ), .ZN(\seg1/_14_ ) );
NOR2_X4 \seg1/_42_ ( .A1(\seg1/_00_ ), .A2(\seg1/_01_ ), .ZN(\seg1/_15_ ) );
INV_X32 \seg1/_43_ ( .A(\seg1/_02_ ), .ZN(\seg1/_16_ ) );
NOR2_X4 \seg1/_44_ ( .A1(\seg1/_16_ ), .A2(\seg1/_03_ ), .ZN(\seg1/_17_ ) );
AOI21_X4 \seg1/_45_ ( .A(\seg1/_14_ ), .B1(\seg1/_15_ ), .B2(\seg1/_17_ ), .ZN(\seg1/_18_ ) );
AND2_X4 \seg1/_46_ ( .A1(\seg1/_00_ ), .A2(\seg1/_01_ ), .ZN(\seg1/_19_ ) );
AND3_X2 \seg1/_47_ ( .A1(\seg1/_19_ ), .A2(\seg1/_03_ ), .A3(\seg1/_16_ ), .ZN(\seg1/_20_ ) );
NOR2_X4 \seg1/_48_ ( .A1(\seg1/_03_ ), .A2(\seg1/_02_ ), .ZN(\seg1/_21_ ) );
AND2_X1 \seg1/_49_ ( .A1(\seg1/_15_ ), .A2(\seg1/_21_ ), .ZN(\seg1/_22_ ) );
NOR2_X2 \seg1/_50_ ( .A1(\seg1/_20_ ), .A2(\seg1/_22_ ), .ZN(\seg1/_23_ ) );
INV_X1 \seg1/_51_ ( .A(\seg1/_21_ ), .ZN(\seg1/_24_ ) );
INV_X1 \seg1/_52_ ( .A(\seg1/_12_ ), .ZN(\seg1/_25_ ) );
OAI211_X2 \seg1/_53_ ( .A(\seg1/_18_ ), .B(\seg1/_23_ ), .C1(\seg1/_24_ ), .C2(\seg1/_25_ ), .ZN(\seg1/_04_ ) );
INV_X16 \seg1/_54_ ( .A(\seg1/_01_ ), .ZN(\seg1/_26_ ) );
NOR2_X4 \seg1/_55_ ( .A1(\seg1/_26_ ), .A2(\seg1/_00_ ), .ZN(\seg1/_27_ ) );
OAI21_X1 \seg1/_56_ ( .A(\seg1/_17_ ), .B1(\seg1/_12_ ), .B2(\seg1/_27_ ), .ZN(\seg1/_28_ ) );
NAND2_X1 \seg1/_57_ ( .A1(\seg1/_25_ ), .A2(\seg1/_13_ ), .ZN(\seg1/_29_ ) );
NAND3_X1 \seg1/_58_ ( .A1(\seg1/_23_ ), .A2(\seg1/_28_ ), .A3(\seg1/_29_ ), .ZN(\seg1/_05_ ) );
OAI21_X1 \seg1/_59_ ( .A(\seg1/_29_ ), .B1(\seg1/_00_ ), .B2(\seg1/_24_ ), .ZN(\seg1/_06_ ) );
INV_X1 \seg1/_60_ ( .A(\seg1/_17_ ), .ZN(\seg1/_30_ ) );
OR3_X2 \seg1/_61_ ( .A1(\seg1/_30_ ), .A2(\seg1/_12_ ), .A3(\seg1/_27_ ), .ZN(\seg1/_31_ ) );
NAND3_X1 \seg1/_62_ ( .A1(\seg1/_27_ ), .A2(\seg1/_03_ ), .A3(\seg1/_16_ ), .ZN(\seg1/_32_ ) );
NAND2_X1 \seg1/_63_ ( .A1(\seg1/_19_ ), .A2(\seg1/_13_ ), .ZN(\seg1/_33_ ) );
NAND2_X1 \seg1/_64_ ( .A1(\seg1/_21_ ), .A2(\seg1/_26_ ), .ZN(\seg1/_34_ ) );
NAND4_X1 \seg1/_65_ ( .A1(\seg1/_31_ ), .A2(\seg1/_32_ ), .A3(\seg1/_33_ ), .A4(\seg1/_34_ ), .ZN(\seg1/_07_ ) );
OAI22_X1 \seg1/_66_ ( .A1(\seg1/_25_ ), .A2(\seg1/_02_ ), .B1(\seg1/_03_ ), .B2(\seg1/_27_ ), .ZN(\seg1/_08_ ) );
AOI22_X1 \seg1/_67_ ( .A1(\seg1/_12_ ), .A2(\seg1/_13_ ), .B1(\seg1/_15_ ), .B2(\seg1/_21_ ), .ZN(\seg1/_35_ ) );
NAND2_X1 \seg1/_68_ ( .A1(\seg1/_17_ ), .A2(\seg1/_19_ ), .ZN(\seg1/_36_ ) );
OAI211_X2 \seg1/_69_ ( .A(\seg1/_35_ ), .B(\seg1/_36_ ), .C1(\seg1/_15_ ), .C2(\seg1/_24_ ), .ZN(\seg1/_09_ ) );
NAND2_X1 \seg1/_70_ ( .A1(\seg1/_13_ ), .A2(\seg1/_15_ ), .ZN(\seg1/_37_ ) );
NAND3_X1 \seg1/_71_ ( .A1(\seg1/_36_ ), .A2(\seg1/_34_ ), .A3(\seg1/_37_ ), .ZN(\seg1/_10_ ) );
BUF_X1 \seg1/_72_ ( .A(\ps2_value[7] ), .Z(\seg1/_03_ ) );
BUF_X1 \seg1/_73_ ( .A(\ps2_value[6] ), .Z(\seg1/_02_ ) );
BUF_X1 \seg1/_74_ ( .A(\ps2_value[4] ), .Z(\seg1/_00_ ) );
BUF_X1 \seg1/_75_ ( .A(\ps2_value[5] ), .Z(\seg1/_01_ ) );
BUF_X1 \seg1/_76_ ( .A(\seg1/_04_ ), .Z(\value_seg[7] ) );
BUF_X1 \seg1/_77_ ( .A(\seg1/_05_ ), .Z(\value_seg[8] ) );
BUF_X1 \seg1/_78_ ( .A(\seg1/_06_ ), .Z(\value_seg[9] ) );
BUF_X1 \seg1/_79_ ( .A(\seg1/_07_ ), .Z(\value_seg[10] ) );
BUF_X1 \seg1/_80_ ( .A(\seg1/_08_ ), .Z(\value_seg[11] ) );
BUF_X1 \seg1/_81_ ( .A(\seg1/_09_ ), .Z(\value_seg[12] ) );
BUF_X1 \seg1/_82_ ( .A(\seg1/_10_ ), .Z(\value_seg[13] ) );
INV_X16 \seg2/_38_ ( .A(\seg2/_00_ ), .ZN(\seg2/_11_ ) );
NOR2_X4 \seg2/_39_ ( .A1(\seg2/_11_ ), .A2(\seg2/_01_ ), .ZN(\seg2/_12_ ) );
AND2_X4 \seg2/_40_ ( .A1(\seg2/_03_ ), .A2(\seg2/_02_ ), .ZN(\seg2/_13_ ) );
AND2_X4 \seg2/_41_ ( .A1(\seg2/_12_ ), .A2(\seg2/_13_ ), .ZN(\seg2/_14_ ) );
NOR2_X4 \seg2/_42_ ( .A1(\seg2/_00_ ), .A2(\seg2/_01_ ), .ZN(\seg2/_15_ ) );
INV_X32 \seg2/_43_ ( .A(\seg2/_02_ ), .ZN(\seg2/_16_ ) );
NOR2_X4 \seg2/_44_ ( .A1(\seg2/_16_ ), .A2(\seg2/_03_ ), .ZN(\seg2/_17_ ) );
AOI21_X4 \seg2/_45_ ( .A(\seg2/_14_ ), .B1(\seg2/_15_ ), .B2(\seg2/_17_ ), .ZN(\seg2/_18_ ) );
AND2_X4 \seg2/_46_ ( .A1(\seg2/_00_ ), .A2(\seg2/_01_ ), .ZN(\seg2/_19_ ) );
AND3_X2 \seg2/_47_ ( .A1(\seg2/_19_ ), .A2(\seg2/_03_ ), .A3(\seg2/_16_ ), .ZN(\seg2/_20_ ) );
NOR2_X4 \seg2/_48_ ( .A1(\seg2/_03_ ), .A2(\seg2/_02_ ), .ZN(\seg2/_21_ ) );
AND2_X1 \seg2/_49_ ( .A1(\seg2/_15_ ), .A2(\seg2/_21_ ), .ZN(\seg2/_22_ ) );
NOR2_X2 \seg2/_50_ ( .A1(\seg2/_20_ ), .A2(\seg2/_22_ ), .ZN(\seg2/_23_ ) );
INV_X1 \seg2/_51_ ( .A(\seg2/_21_ ), .ZN(\seg2/_24_ ) );
INV_X1 \seg2/_52_ ( .A(\seg2/_12_ ), .ZN(\seg2/_25_ ) );
OAI211_X2 \seg2/_53_ ( .A(\seg2/_18_ ), .B(\seg2/_23_ ), .C1(\seg2/_24_ ), .C2(\seg2/_25_ ), .ZN(\seg2/_04_ ) );
INV_X16 \seg2/_54_ ( .A(\seg2/_01_ ), .ZN(\seg2/_26_ ) );
NOR2_X4 \seg2/_55_ ( .A1(\seg2/_26_ ), .A2(\seg2/_00_ ), .ZN(\seg2/_27_ ) );
OAI21_X1 \seg2/_56_ ( .A(\seg2/_17_ ), .B1(\seg2/_12_ ), .B2(\seg2/_27_ ), .ZN(\seg2/_28_ ) );
NAND2_X1 \seg2/_57_ ( .A1(\seg2/_25_ ), .A2(\seg2/_13_ ), .ZN(\seg2/_29_ ) );
NAND3_X1 \seg2/_58_ ( .A1(\seg2/_23_ ), .A2(\seg2/_28_ ), .A3(\seg2/_29_ ), .ZN(\seg2/_05_ ) );
OAI21_X1 \seg2/_59_ ( .A(\seg2/_29_ ), .B1(\seg2/_00_ ), .B2(\seg2/_24_ ), .ZN(\seg2/_06_ ) );
INV_X1 \seg2/_60_ ( .A(\seg2/_17_ ), .ZN(\seg2/_30_ ) );
OR3_X2 \seg2/_61_ ( .A1(\seg2/_30_ ), .A2(\seg2/_12_ ), .A3(\seg2/_27_ ), .ZN(\seg2/_31_ ) );
NAND3_X1 \seg2/_62_ ( .A1(\seg2/_27_ ), .A2(\seg2/_03_ ), .A3(\seg2/_16_ ), .ZN(\seg2/_32_ ) );
NAND2_X1 \seg2/_63_ ( .A1(\seg2/_19_ ), .A2(\seg2/_13_ ), .ZN(\seg2/_33_ ) );
NAND2_X1 \seg2/_64_ ( .A1(\seg2/_21_ ), .A2(\seg2/_26_ ), .ZN(\seg2/_34_ ) );
NAND4_X1 \seg2/_65_ ( .A1(\seg2/_31_ ), .A2(\seg2/_32_ ), .A3(\seg2/_33_ ), .A4(\seg2/_34_ ), .ZN(\seg2/_07_ ) );
OAI22_X1 \seg2/_66_ ( .A1(\seg2/_25_ ), .A2(\seg2/_02_ ), .B1(\seg2/_03_ ), .B2(\seg2/_27_ ), .ZN(\seg2/_08_ ) );
AOI22_X1 \seg2/_67_ ( .A1(\seg2/_12_ ), .A2(\seg2/_13_ ), .B1(\seg2/_15_ ), .B2(\seg2/_21_ ), .ZN(\seg2/_35_ ) );
NAND2_X1 \seg2/_68_ ( .A1(\seg2/_17_ ), .A2(\seg2/_19_ ), .ZN(\seg2/_36_ ) );
OAI211_X2 \seg2/_69_ ( .A(\seg2/_35_ ), .B(\seg2/_36_ ), .C1(\seg2/_15_ ), .C2(\seg2/_24_ ), .ZN(\seg2/_09_ ) );
NAND2_X1 \seg2/_70_ ( .A1(\seg2/_13_ ), .A2(\seg2/_15_ ), .ZN(\seg2/_37_ ) );
NAND3_X1 \seg2/_71_ ( .A1(\seg2/_36_ ), .A2(\seg2/_34_ ), .A3(\seg2/_37_ ), .ZN(\seg2/_10_ ) );
BUF_X1 \seg2/_72_ ( .A(\ps2_value[11] ), .Z(\seg2/_03_ ) );
BUF_X1 \seg2/_73_ ( .A(\ps2_value[10] ), .Z(\seg2/_02_ ) );
BUF_X1 \seg2/_74_ ( .A(\ps2_value[8] ), .Z(\seg2/_00_ ) );
BUF_X1 \seg2/_75_ ( .A(\ps2_value[9] ), .Z(\seg2/_01_ ) );
BUF_X1 \seg2/_76_ ( .A(\seg2/_04_ ), .Z(\value_seg[14] ) );
BUF_X1 \seg2/_77_ ( .A(\seg2/_05_ ), .Z(\value_seg[15] ) );
BUF_X1 \seg2/_78_ ( .A(\seg2/_06_ ), .Z(\value_seg[16] ) );
BUF_X1 \seg2/_79_ ( .A(\seg2/_07_ ), .Z(\value_seg[17] ) );
BUF_X1 \seg2/_80_ ( .A(\seg2/_08_ ), .Z(\value_seg[18] ) );
BUF_X1 \seg2/_81_ ( .A(\seg2/_09_ ), .Z(\value_seg[19] ) );
BUF_X1 \seg2/_82_ ( .A(\seg2/_10_ ), .Z(\value_seg[20] ) );
INV_X16 \seg3/_38_ ( .A(\seg3/_00_ ), .ZN(\seg3/_11_ ) );
NOR2_X4 \seg3/_39_ ( .A1(\seg3/_11_ ), .A2(\seg3/_01_ ), .ZN(\seg3/_12_ ) );
AND2_X4 \seg3/_40_ ( .A1(\seg3/_03_ ), .A2(\seg3/_02_ ), .ZN(\seg3/_13_ ) );
AND2_X4 \seg3/_41_ ( .A1(\seg3/_12_ ), .A2(\seg3/_13_ ), .ZN(\seg3/_14_ ) );
NOR2_X4 \seg3/_42_ ( .A1(\seg3/_00_ ), .A2(\seg3/_01_ ), .ZN(\seg3/_15_ ) );
INV_X32 \seg3/_43_ ( .A(\seg3/_02_ ), .ZN(\seg3/_16_ ) );
NOR2_X4 \seg3/_44_ ( .A1(\seg3/_16_ ), .A2(\seg3/_03_ ), .ZN(\seg3/_17_ ) );
AOI21_X4 \seg3/_45_ ( .A(\seg3/_14_ ), .B1(\seg3/_15_ ), .B2(\seg3/_17_ ), .ZN(\seg3/_18_ ) );
AND2_X4 \seg3/_46_ ( .A1(\seg3/_00_ ), .A2(\seg3/_01_ ), .ZN(\seg3/_19_ ) );
AND3_X2 \seg3/_47_ ( .A1(\seg3/_19_ ), .A2(\seg3/_03_ ), .A3(\seg3/_16_ ), .ZN(\seg3/_20_ ) );
NOR2_X4 \seg3/_48_ ( .A1(\seg3/_03_ ), .A2(\seg3/_02_ ), .ZN(\seg3/_21_ ) );
AND2_X1 \seg3/_49_ ( .A1(\seg3/_15_ ), .A2(\seg3/_21_ ), .ZN(\seg3/_22_ ) );
NOR2_X2 \seg3/_50_ ( .A1(\seg3/_20_ ), .A2(\seg3/_22_ ), .ZN(\seg3/_23_ ) );
INV_X1 \seg3/_51_ ( .A(\seg3/_21_ ), .ZN(\seg3/_24_ ) );
INV_X1 \seg3/_52_ ( .A(\seg3/_12_ ), .ZN(\seg3/_25_ ) );
OAI211_X2 \seg3/_53_ ( .A(\seg3/_18_ ), .B(\seg3/_23_ ), .C1(\seg3/_24_ ), .C2(\seg3/_25_ ), .ZN(\seg3/_04_ ) );
INV_X16 \seg3/_54_ ( .A(\seg3/_01_ ), .ZN(\seg3/_26_ ) );
NOR2_X4 \seg3/_55_ ( .A1(\seg3/_26_ ), .A2(\seg3/_00_ ), .ZN(\seg3/_27_ ) );
OAI21_X1 \seg3/_56_ ( .A(\seg3/_17_ ), .B1(\seg3/_12_ ), .B2(\seg3/_27_ ), .ZN(\seg3/_28_ ) );
NAND2_X1 \seg3/_57_ ( .A1(\seg3/_25_ ), .A2(\seg3/_13_ ), .ZN(\seg3/_29_ ) );
NAND3_X1 \seg3/_58_ ( .A1(\seg3/_23_ ), .A2(\seg3/_28_ ), .A3(\seg3/_29_ ), .ZN(\seg3/_05_ ) );
OAI21_X1 \seg3/_59_ ( .A(\seg3/_29_ ), .B1(\seg3/_00_ ), .B2(\seg3/_24_ ), .ZN(\seg3/_06_ ) );
INV_X1 \seg3/_60_ ( .A(\seg3/_17_ ), .ZN(\seg3/_30_ ) );
OR3_X2 \seg3/_61_ ( .A1(\seg3/_30_ ), .A2(\seg3/_12_ ), .A3(\seg3/_27_ ), .ZN(\seg3/_31_ ) );
NAND3_X1 \seg3/_62_ ( .A1(\seg3/_27_ ), .A2(\seg3/_03_ ), .A3(\seg3/_16_ ), .ZN(\seg3/_32_ ) );
NAND2_X1 \seg3/_63_ ( .A1(\seg3/_19_ ), .A2(\seg3/_13_ ), .ZN(\seg3/_33_ ) );
NAND2_X1 \seg3/_64_ ( .A1(\seg3/_21_ ), .A2(\seg3/_26_ ), .ZN(\seg3/_34_ ) );
NAND4_X1 \seg3/_65_ ( .A1(\seg3/_31_ ), .A2(\seg3/_32_ ), .A3(\seg3/_33_ ), .A4(\seg3/_34_ ), .ZN(\seg3/_07_ ) );
OAI22_X1 \seg3/_66_ ( .A1(\seg3/_25_ ), .A2(\seg3/_02_ ), .B1(\seg3/_03_ ), .B2(\seg3/_27_ ), .ZN(\seg3/_08_ ) );
AOI22_X1 \seg3/_67_ ( .A1(\seg3/_12_ ), .A2(\seg3/_13_ ), .B1(\seg3/_15_ ), .B2(\seg3/_21_ ), .ZN(\seg3/_35_ ) );
NAND2_X1 \seg3/_68_ ( .A1(\seg3/_17_ ), .A2(\seg3/_19_ ), .ZN(\seg3/_36_ ) );
OAI211_X2 \seg3/_69_ ( .A(\seg3/_35_ ), .B(\seg3/_36_ ), .C1(\seg3/_15_ ), .C2(\seg3/_24_ ), .ZN(\seg3/_09_ ) );
NAND2_X1 \seg3/_70_ ( .A1(\seg3/_13_ ), .A2(\seg3/_15_ ), .ZN(\seg3/_37_ ) );
NAND3_X1 \seg3/_71_ ( .A1(\seg3/_36_ ), .A2(\seg3/_34_ ), .A3(\seg3/_37_ ), .ZN(\seg3/_10_ ) );
BUF_X1 \seg3/_72_ ( .A(\ps2_value[15] ), .Z(\seg3/_03_ ) );
BUF_X1 \seg3/_73_ ( .A(\ps2_value[14] ), .Z(\seg3/_02_ ) );
BUF_X1 \seg3/_74_ ( .A(\ps2_value[12] ), .Z(\seg3/_00_ ) );
BUF_X1 \seg3/_75_ ( .A(\ps2_value[13] ), .Z(\seg3/_01_ ) );
BUF_X1 \seg3/_76_ ( .A(\seg3/_04_ ), .Z(\value_seg[21] ) );
BUF_X1 \seg3/_77_ ( .A(\seg3/_05_ ), .Z(\value_seg[22] ) );
BUF_X1 \seg3/_78_ ( .A(\seg3/_06_ ), .Z(\value_seg[23] ) );
BUF_X1 \seg3/_79_ ( .A(\seg3/_07_ ), .Z(\value_seg[24] ) );
BUF_X1 \seg3/_80_ ( .A(\seg3/_08_ ), .Z(\value_seg[25] ) );
BUF_X1 \seg3/_81_ ( .A(\seg3/_09_ ), .Z(\value_seg[26] ) );
BUF_X1 \seg3/_82_ ( .A(\seg3/_10_ ), .Z(\value_seg[27] ) );
INV_X16 \seg4/_38_ ( .A(\seg4/_00_ ), .ZN(\seg4/_11_ ) );
NOR2_X4 \seg4/_39_ ( .A1(\seg4/_11_ ), .A2(\seg4/_01_ ), .ZN(\seg4/_12_ ) );
AND2_X4 \seg4/_40_ ( .A1(\seg4/_03_ ), .A2(\seg4/_02_ ), .ZN(\seg4/_13_ ) );
AND2_X4 \seg4/_41_ ( .A1(\seg4/_12_ ), .A2(\seg4/_13_ ), .ZN(\seg4/_14_ ) );
NOR2_X4 \seg4/_42_ ( .A1(\seg4/_00_ ), .A2(\seg4/_01_ ), .ZN(\seg4/_15_ ) );
INV_X32 \seg4/_43_ ( .A(\seg4/_02_ ), .ZN(\seg4/_16_ ) );
NOR2_X4 \seg4/_44_ ( .A1(\seg4/_16_ ), .A2(\seg4/_03_ ), .ZN(\seg4/_17_ ) );
AOI21_X4 \seg4/_45_ ( .A(\seg4/_14_ ), .B1(\seg4/_15_ ), .B2(\seg4/_17_ ), .ZN(\seg4/_18_ ) );
AND2_X4 \seg4/_46_ ( .A1(\seg4/_00_ ), .A2(\seg4/_01_ ), .ZN(\seg4/_19_ ) );
AND3_X2 \seg4/_47_ ( .A1(\seg4/_19_ ), .A2(\seg4/_03_ ), .A3(\seg4/_16_ ), .ZN(\seg4/_20_ ) );
NOR2_X4 \seg4/_48_ ( .A1(\seg4/_03_ ), .A2(\seg4/_02_ ), .ZN(\seg4/_21_ ) );
AND2_X1 \seg4/_49_ ( .A1(\seg4/_15_ ), .A2(\seg4/_21_ ), .ZN(\seg4/_22_ ) );
NOR2_X2 \seg4/_50_ ( .A1(\seg4/_20_ ), .A2(\seg4/_22_ ), .ZN(\seg4/_23_ ) );
INV_X1 \seg4/_51_ ( .A(\seg4/_21_ ), .ZN(\seg4/_24_ ) );
INV_X1 \seg4/_52_ ( .A(\seg4/_12_ ), .ZN(\seg4/_25_ ) );
OAI211_X2 \seg4/_53_ ( .A(\seg4/_18_ ), .B(\seg4/_23_ ), .C1(\seg4/_24_ ), .C2(\seg4/_25_ ), .ZN(\seg4/_04_ ) );
INV_X16 \seg4/_54_ ( .A(\seg4/_01_ ), .ZN(\seg4/_26_ ) );
NOR2_X4 \seg4/_55_ ( .A1(\seg4/_26_ ), .A2(\seg4/_00_ ), .ZN(\seg4/_27_ ) );
OAI21_X1 \seg4/_56_ ( .A(\seg4/_17_ ), .B1(\seg4/_12_ ), .B2(\seg4/_27_ ), .ZN(\seg4/_28_ ) );
NAND2_X1 \seg4/_57_ ( .A1(\seg4/_25_ ), .A2(\seg4/_13_ ), .ZN(\seg4/_29_ ) );
NAND3_X1 \seg4/_58_ ( .A1(\seg4/_23_ ), .A2(\seg4/_28_ ), .A3(\seg4/_29_ ), .ZN(\seg4/_05_ ) );
OAI21_X1 \seg4/_59_ ( .A(\seg4/_29_ ), .B1(\seg4/_00_ ), .B2(\seg4/_24_ ), .ZN(\seg4/_06_ ) );
INV_X1 \seg4/_60_ ( .A(\seg4/_17_ ), .ZN(\seg4/_30_ ) );
OR3_X2 \seg4/_61_ ( .A1(\seg4/_30_ ), .A2(\seg4/_12_ ), .A3(\seg4/_27_ ), .ZN(\seg4/_31_ ) );
NAND3_X1 \seg4/_62_ ( .A1(\seg4/_27_ ), .A2(\seg4/_03_ ), .A3(\seg4/_16_ ), .ZN(\seg4/_32_ ) );
NAND2_X1 \seg4/_63_ ( .A1(\seg4/_19_ ), .A2(\seg4/_13_ ), .ZN(\seg4/_33_ ) );
NAND2_X1 \seg4/_64_ ( .A1(\seg4/_21_ ), .A2(\seg4/_26_ ), .ZN(\seg4/_34_ ) );
NAND4_X1 \seg4/_65_ ( .A1(\seg4/_31_ ), .A2(\seg4/_32_ ), .A3(\seg4/_33_ ), .A4(\seg4/_34_ ), .ZN(\seg4/_07_ ) );
OAI22_X1 \seg4/_66_ ( .A1(\seg4/_25_ ), .A2(\seg4/_02_ ), .B1(\seg4/_03_ ), .B2(\seg4/_27_ ), .ZN(\seg4/_08_ ) );
AOI22_X1 \seg4/_67_ ( .A1(\seg4/_12_ ), .A2(\seg4/_13_ ), .B1(\seg4/_15_ ), .B2(\seg4/_21_ ), .ZN(\seg4/_35_ ) );
NAND2_X1 \seg4/_68_ ( .A1(\seg4/_17_ ), .A2(\seg4/_19_ ), .ZN(\seg4/_36_ ) );
OAI211_X2 \seg4/_69_ ( .A(\seg4/_35_ ), .B(\seg4/_36_ ), .C1(\seg4/_15_ ), .C2(\seg4/_24_ ), .ZN(\seg4/_09_ ) );
NAND2_X1 \seg4/_70_ ( .A1(\seg4/_13_ ), .A2(\seg4/_15_ ), .ZN(\seg4/_37_ ) );
NAND3_X1 \seg4/_71_ ( .A1(\seg4/_36_ ), .A2(\seg4/_34_ ), .A3(\seg4/_37_ ), .ZN(\seg4/_10_ ) );
BUF_X1 \seg4/_72_ ( .A(\count[3] ), .Z(\seg4/_03_ ) );
BUF_X1 \seg4/_73_ ( .A(\count[2] ), .Z(\seg4/_02_ ) );
BUF_X1 \seg4/_74_ ( .A(\count[0] ), .Z(\seg4/_00_ ) );
BUF_X1 \seg4/_75_ ( .A(\count[1] ), .Z(\seg4/_01_ ) );
BUF_X1 \seg4/_76_ ( .A(\seg4/_04_ ), .Z(\value_seg[28] ) );
BUF_X1 \seg4/_77_ ( .A(\seg4/_05_ ), .Z(\value_seg[29] ) );
BUF_X1 \seg4/_78_ ( .A(\seg4/_06_ ), .Z(\value_seg[30] ) );
BUF_X1 \seg4/_79_ ( .A(\seg4/_07_ ), .Z(\value_seg[31] ) );
BUF_X1 \seg4/_80_ ( .A(\seg4/_08_ ), .Z(\value_seg[32] ) );
BUF_X1 \seg4/_81_ ( .A(\seg4/_09_ ), .Z(\value_seg[33] ) );
BUF_X1 \seg4/_82_ ( .A(\seg4/_10_ ), .Z(\value_seg[34] ) );
INV_X16 \seg5/_38_ ( .A(\seg5/_00_ ), .ZN(\seg5/_11_ ) );
NOR2_X4 \seg5/_39_ ( .A1(\seg5/_11_ ), .A2(\seg5/_01_ ), .ZN(\seg5/_12_ ) );
AND2_X4 \seg5/_40_ ( .A1(\seg5/_03_ ), .A2(\seg5/_02_ ), .ZN(\seg5/_13_ ) );
AND2_X4 \seg5/_41_ ( .A1(\seg5/_12_ ), .A2(\seg5/_13_ ), .ZN(\seg5/_14_ ) );
NOR2_X4 \seg5/_42_ ( .A1(\seg5/_00_ ), .A2(\seg5/_01_ ), .ZN(\seg5/_15_ ) );
INV_X32 \seg5/_43_ ( .A(\seg5/_02_ ), .ZN(\seg5/_16_ ) );
NOR2_X4 \seg5/_44_ ( .A1(\seg5/_16_ ), .A2(\seg5/_03_ ), .ZN(\seg5/_17_ ) );
AOI21_X4 \seg5/_45_ ( .A(\seg5/_14_ ), .B1(\seg5/_15_ ), .B2(\seg5/_17_ ), .ZN(\seg5/_18_ ) );
AND2_X4 \seg5/_46_ ( .A1(\seg5/_00_ ), .A2(\seg5/_01_ ), .ZN(\seg5/_19_ ) );
AND3_X2 \seg5/_47_ ( .A1(\seg5/_19_ ), .A2(\seg5/_03_ ), .A3(\seg5/_16_ ), .ZN(\seg5/_20_ ) );
NOR2_X4 \seg5/_48_ ( .A1(\seg5/_03_ ), .A2(\seg5/_02_ ), .ZN(\seg5/_21_ ) );
AND2_X1 \seg5/_49_ ( .A1(\seg5/_15_ ), .A2(\seg5/_21_ ), .ZN(\seg5/_22_ ) );
NOR2_X2 \seg5/_50_ ( .A1(\seg5/_20_ ), .A2(\seg5/_22_ ), .ZN(\seg5/_23_ ) );
INV_X1 \seg5/_51_ ( .A(\seg5/_21_ ), .ZN(\seg5/_24_ ) );
INV_X1 \seg5/_52_ ( .A(\seg5/_12_ ), .ZN(\seg5/_25_ ) );
OAI211_X2 \seg5/_53_ ( .A(\seg5/_18_ ), .B(\seg5/_23_ ), .C1(\seg5/_24_ ), .C2(\seg5/_25_ ), .ZN(\seg5/_04_ ) );
INV_X16 \seg5/_54_ ( .A(\seg5/_01_ ), .ZN(\seg5/_26_ ) );
NOR2_X4 \seg5/_55_ ( .A1(\seg5/_26_ ), .A2(\seg5/_00_ ), .ZN(\seg5/_27_ ) );
OAI21_X1 \seg5/_56_ ( .A(\seg5/_17_ ), .B1(\seg5/_12_ ), .B2(\seg5/_27_ ), .ZN(\seg5/_28_ ) );
NAND2_X1 \seg5/_57_ ( .A1(\seg5/_25_ ), .A2(\seg5/_13_ ), .ZN(\seg5/_29_ ) );
NAND3_X1 \seg5/_58_ ( .A1(\seg5/_23_ ), .A2(\seg5/_28_ ), .A3(\seg5/_29_ ), .ZN(\seg5/_05_ ) );
OAI21_X1 \seg5/_59_ ( .A(\seg5/_29_ ), .B1(\seg5/_00_ ), .B2(\seg5/_24_ ), .ZN(\seg5/_06_ ) );
INV_X1 \seg5/_60_ ( .A(\seg5/_17_ ), .ZN(\seg5/_30_ ) );
OR3_X2 \seg5/_61_ ( .A1(\seg5/_30_ ), .A2(\seg5/_12_ ), .A3(\seg5/_27_ ), .ZN(\seg5/_31_ ) );
NAND3_X1 \seg5/_62_ ( .A1(\seg5/_27_ ), .A2(\seg5/_03_ ), .A3(\seg5/_16_ ), .ZN(\seg5/_32_ ) );
NAND2_X1 \seg5/_63_ ( .A1(\seg5/_19_ ), .A2(\seg5/_13_ ), .ZN(\seg5/_33_ ) );
NAND2_X1 \seg5/_64_ ( .A1(\seg5/_21_ ), .A2(\seg5/_26_ ), .ZN(\seg5/_34_ ) );
NAND4_X1 \seg5/_65_ ( .A1(\seg5/_31_ ), .A2(\seg5/_32_ ), .A3(\seg5/_33_ ), .A4(\seg5/_34_ ), .ZN(\seg5/_07_ ) );
OAI22_X1 \seg5/_66_ ( .A1(\seg5/_25_ ), .A2(\seg5/_02_ ), .B1(\seg5/_03_ ), .B2(\seg5/_27_ ), .ZN(\seg5/_08_ ) );
AOI22_X1 \seg5/_67_ ( .A1(\seg5/_12_ ), .A2(\seg5/_13_ ), .B1(\seg5/_15_ ), .B2(\seg5/_21_ ), .ZN(\seg5/_35_ ) );
NAND2_X1 \seg5/_68_ ( .A1(\seg5/_17_ ), .A2(\seg5/_19_ ), .ZN(\seg5/_36_ ) );
OAI211_X2 \seg5/_69_ ( .A(\seg5/_35_ ), .B(\seg5/_36_ ), .C1(\seg5/_15_ ), .C2(\seg5/_24_ ), .ZN(\seg5/_09_ ) );
NAND2_X1 \seg5/_70_ ( .A1(\seg5/_13_ ), .A2(\seg5/_15_ ), .ZN(\seg5/_37_ ) );
NAND3_X1 \seg5/_71_ ( .A1(\seg5/_36_ ), .A2(\seg5/_34_ ), .A3(\seg5/_37_ ), .ZN(\seg5/_10_ ) );
BUF_X1 \seg5/_72_ ( .A(\count[7] ), .Z(\seg5/_03_ ) );
BUF_X1 \seg5/_73_ ( .A(\count[6] ), .Z(\seg5/_02_ ) );
BUF_X1 \seg5/_74_ ( .A(\count[4] ), .Z(\seg5/_00_ ) );
BUF_X1 \seg5/_75_ ( .A(\count[5] ), .Z(\seg5/_01_ ) );
BUF_X1 \seg5/_76_ ( .A(\seg5/_04_ ), .Z(\value_seg[35] ) );
BUF_X1 \seg5/_77_ ( .A(\seg5/_05_ ), .Z(\value_seg[36] ) );
BUF_X1 \seg5/_78_ ( .A(\seg5/_06_ ), .Z(\value_seg[37] ) );
BUF_X1 \seg5/_79_ ( .A(\seg5/_07_ ), .Z(\value_seg[38] ) );
BUF_X1 \seg5/_80_ ( .A(\seg5/_08_ ), .Z(\value_seg[39] ) );
BUF_X1 \seg5/_81_ ( .A(\seg5/_09_ ), .Z(\value_seg[40] ) );
BUF_X1 \seg5/_82_ ( .A(\seg5/_10_ ), .Z(\value_seg[41] ) );

endmodule
