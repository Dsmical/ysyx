//Generate the verilog at 2024-03-17T14:44:03
module gcd (
clk,
req_rdy,
req_val,
reset,
resp_rdy,
resp_val,
req_msg,
resp_msg
);

input clk ;
output req_rdy ;
input req_val ;
input reset ;
input resp_rdy ;
output resp_val ;
input [31:0] req_msg ;
output [15:0] resp_msg ;

wire \ctrl$a_mux_sel[0] ;
wire \ctrl$a_mux_sel[1] ;
wire ctrl$a_reg_en ;
wire ctrl$b_mux_sel ;
wire ctrl$b_reg_en ;
wire ctrl$is_a_lt_b ;
wire ctrl$is_b_zero ;
wire \ctrl/_00_ ;
wire \ctrl/_01_ ;
wire \ctrl/_02_ ;
wire \ctrl/_03_ ;
wire \ctrl/_04_ ;
wire \ctrl/_05_ ;
wire \ctrl/_06_ ;
wire \ctrl/_07_ ;
wire \ctrl/_08_ ;
wire \ctrl/_09_ ;
wire \ctrl/_10_ ;
wire \ctrl/_11_ ;
wire \ctrl/_12_ ;
wire \ctrl/_13_ ;
wire \ctrl/_14_ ;
wire \ctrl/_15_ ;
wire \ctrl/_16_ ;
wire \ctrl/_17_ ;
wire \ctrl/_18_ ;
wire \ctrl/_19_ ;
wire \ctrl/curr_state__0[0] ;
wire \ctrl/curr_state__0[1] ;
wire \ctrl/next_state__0[0] ;
wire \ctrl/next_state__0[1] ;
wire req_rdy ;
wire resp_val ;
wire req_val ;
wire resp_rdy ;
wire \ctrl/state/_00_ ;
wire \ctrl/state/_01_ ;
wire \ctrl/state/_02_ ;
wire \ctrl/state/_03_ ;
wire \ctrl/state/_04_ ;
wire \ctrl/state/_05_ ;
wire \ctrl/state/_06_ ;
wire \ctrl/state/_07_ ;
wire \ctrl/state/_08_ ;
wire \ctrl/state/_09_ ;
wire \ctrl/state/_10_ ;
wire reset ;
wire clk ;
wire \dpath/a_lt_b$in0[0] ;
wire \dpath/a_lt_b$in0[10] ;
wire \dpath/a_lt_b$in0[11] ;
wire \dpath/a_lt_b$in0[12] ;
wire \dpath/a_lt_b$in0[13] ;
wire \dpath/a_lt_b$in0[14] ;
wire \dpath/a_lt_b$in0[15] ;
wire \dpath/a_lt_b$in0[1] ;
wire \dpath/a_lt_b$in0[2] ;
wire \dpath/a_lt_b$in0[3] ;
wire \dpath/a_lt_b$in0[4] ;
wire \dpath/a_lt_b$in0[5] ;
wire \dpath/a_lt_b$in0[6] ;
wire \dpath/a_lt_b$in0[7] ;
wire \dpath/a_lt_b$in0[8] ;
wire \dpath/a_lt_b$in0[9] ;
wire \dpath/a_lt_b$in1[0] ;
wire \dpath/a_lt_b$in1[10] ;
wire \dpath/a_lt_b$in1[11] ;
wire \dpath/a_lt_b$in1[12] ;
wire \dpath/a_lt_b$in1[13] ;
wire \dpath/a_lt_b$in1[14] ;
wire \dpath/a_lt_b$in1[15] ;
wire \dpath/a_lt_b$in1[1] ;
wire \dpath/a_lt_b$in1[2] ;
wire \dpath/a_lt_b$in1[3] ;
wire \dpath/a_lt_b$in1[4] ;
wire \dpath/a_lt_b$in1[5] ;
wire \dpath/a_lt_b$in1[6] ;
wire \dpath/a_lt_b$in1[7] ;
wire \dpath/a_lt_b$in1[8] ;
wire \dpath/a_lt_b$in1[9] ;
wire \dpath/a_mux$out[0] ;
wire \dpath/a_mux$out[10] ;
wire \dpath/a_mux$out[11] ;
wire \dpath/a_mux$out[12] ;
wire \dpath/a_mux$out[13] ;
wire \dpath/a_mux$out[14] ;
wire \dpath/a_mux$out[15] ;
wire \dpath/a_mux$out[1] ;
wire \dpath/a_mux$out[2] ;
wire \dpath/a_mux$out[3] ;
wire \dpath/a_mux$out[4] ;
wire \dpath/a_mux$out[5] ;
wire \dpath/a_mux$out[6] ;
wire \dpath/a_mux$out[7] ;
wire \dpath/a_mux$out[8] ;
wire \dpath/a_mux$out[9] ;
wire \dpath/b_mux$out[0] ;
wire \dpath/b_mux$out[10] ;
wire \dpath/b_mux$out[11] ;
wire \dpath/b_mux$out[12] ;
wire \dpath/b_mux$out[13] ;
wire \dpath/b_mux$out[14] ;
wire \dpath/b_mux$out[15] ;
wire \dpath/b_mux$out[1] ;
wire \dpath/b_mux$out[2] ;
wire \dpath/b_mux$out[3] ;
wire \dpath/b_mux$out[4] ;
wire \dpath/b_mux$out[5] ;
wire \dpath/b_mux$out[6] ;
wire \dpath/b_mux$out[7] ;
wire \dpath/b_mux$out[8] ;
wire \dpath/b_mux$out[9] ;
wire \dpath/a_lt_b/_000_ ;
wire \dpath/a_lt_b/_001_ ;
wire \dpath/a_lt_b/_002_ ;
wire \dpath/a_lt_b/_003_ ;
wire \dpath/a_lt_b/_004_ ;
wire \dpath/a_lt_b/_005_ ;
wire \dpath/a_lt_b/_006_ ;
wire \dpath/a_lt_b/_007_ ;
wire \dpath/a_lt_b/_008_ ;
wire \dpath/a_lt_b/_009_ ;
wire \dpath/a_lt_b/_010_ ;
wire \dpath/a_lt_b/_011_ ;
wire \dpath/a_lt_b/_012_ ;
wire \dpath/a_lt_b/_013_ ;
wire \dpath/a_lt_b/_014_ ;
wire \dpath/a_lt_b/_015_ ;
wire \dpath/a_lt_b/_016_ ;
wire \dpath/a_lt_b/_017_ ;
wire \dpath/a_lt_b/_018_ ;
wire \dpath/a_lt_b/_019_ ;
wire \dpath/a_lt_b/_020_ ;
wire \dpath/a_lt_b/_021_ ;
wire \dpath/a_lt_b/_022_ ;
wire \dpath/a_lt_b/_023_ ;
wire \dpath/a_lt_b/_024_ ;
wire \dpath/a_lt_b/_025_ ;
wire \dpath/a_lt_b/_026_ ;
wire \dpath/a_lt_b/_027_ ;
wire \dpath/a_lt_b/_028_ ;
wire \dpath/a_lt_b/_029_ ;
wire \dpath/a_lt_b/_030_ ;
wire \dpath/a_lt_b/_031_ ;
wire \dpath/a_lt_b/_032_ ;
wire \dpath/a_lt_b/_033_ ;
wire \dpath/a_lt_b/_034_ ;
wire \dpath/a_lt_b/_035_ ;
wire \dpath/a_lt_b/_036_ ;
wire \dpath/a_lt_b/_037_ ;
wire \dpath/a_lt_b/_038_ ;
wire \dpath/a_lt_b/_039_ ;
wire \dpath/a_lt_b/_040_ ;
wire \dpath/a_lt_b/_041_ ;
wire \dpath/a_lt_b/_042_ ;
wire \dpath/a_lt_b/_043_ ;
wire \dpath/a_lt_b/_044_ ;
wire \dpath/a_lt_b/_045_ ;
wire \dpath/a_lt_b/_046_ ;
wire \dpath/a_lt_b/_047_ ;
wire \dpath/a_lt_b/_048_ ;
wire \dpath/a_lt_b/_049_ ;
wire \dpath/a_lt_b/_050_ ;
wire \dpath/a_lt_b/_051_ ;
wire \dpath/a_lt_b/_052_ ;
wire \dpath/a_lt_b/_053_ ;
wire \dpath/a_lt_b/_054_ ;
wire \dpath/a_lt_b/_055_ ;
wire \dpath/a_lt_b/_056_ ;
wire \dpath/a_lt_b/_057_ ;
wire \dpath/a_lt_b/_058_ ;
wire \dpath/a_lt_b/_059_ ;
wire \dpath/a_lt_b/_060_ ;
wire \dpath/a_lt_b/_061_ ;
wire \dpath/a_lt_b/_062_ ;
wire \dpath/a_lt_b/_063_ ;
wire \dpath/a_lt_b/_064_ ;
wire \dpath/a_lt_b/_065_ ;
wire \dpath/a_lt_b/_066_ ;
wire \dpath/a_lt_b/_067_ ;
wire \dpath/a_lt_b/_068_ ;
wire \dpath/a_lt_b/_069_ ;
wire \dpath/a_lt_b/_070_ ;
wire \dpath/a_lt_b/_071_ ;
wire \dpath/a_lt_b/_072_ ;
wire \dpath/a_lt_b/_073_ ;
wire \dpath/a_lt_b/_074_ ;
wire \dpath/a_lt_b/_075_ ;
wire \dpath/a_lt_b/_076_ ;
wire \dpath/a_lt_b/_077_ ;
wire \dpath/a_lt_b/_078_ ;
wire \dpath/a_lt_b/_079_ ;
wire \dpath/a_lt_b/_080_ ;
wire \dpath/a_lt_b/_081_ ;
wire \dpath/a_lt_b/_082_ ;
wire \dpath/a_lt_b/_083_ ;
wire \dpath/a_lt_b/_084_ ;
wire \dpath/a_lt_b/_085_ ;
wire \dpath/a_lt_b/_086_ ;
wire \dpath/a_lt_b/_087_ ;
wire \dpath/a_lt_b/_088_ ;
wire \dpath/a_lt_b/_089_ ;
wire \dpath/a_lt_b/_090_ ;
wire \dpath/a_lt_b/_091_ ;
wire \dpath/a_lt_b/_092_ ;
wire \dpath/a_lt_b/_093_ ;
wire \dpath/a_lt_b/_094_ ;
wire \dpath/a_lt_b/_095_ ;
wire \dpath/a_lt_b/_096_ ;
wire \dpath/a_lt_b/_097_ ;
wire \dpath/a_lt_b/_098_ ;
wire \dpath/a_lt_b/_099_ ;
wire \dpath/a_lt_b/_100_ ;
wire \dpath/a_lt_b/_101_ ;
wire \dpath/a_lt_b/_102_ ;
wire \dpath/a_lt_b/_103_ ;
wire \dpath/a_lt_b/_104_ ;
wire \dpath/a_lt_b/_105_ ;
wire \dpath/a_lt_b/_106_ ;
wire \dpath/a_lt_b/_107_ ;
wire \dpath/a_lt_b/_108_ ;
wire \dpath/a_mux/_000_ ;
wire \dpath/a_mux/_001_ ;
wire \dpath/a_mux/_002_ ;
wire \dpath/a_mux/_003_ ;
wire \dpath/a_mux/_004_ ;
wire \dpath/a_mux/_005_ ;
wire \dpath/a_mux/_006_ ;
wire \dpath/a_mux/_007_ ;
wire \dpath/a_mux/_008_ ;
wire \dpath/a_mux/_009_ ;
wire \dpath/a_mux/_010_ ;
wire \dpath/a_mux/_011_ ;
wire \dpath/a_mux/_012_ ;
wire \dpath/a_mux/_013_ ;
wire \dpath/a_mux/_014_ ;
wire \dpath/a_mux/_015_ ;
wire \dpath/a_mux/_016_ ;
wire \dpath/a_mux/_017_ ;
wire \dpath/a_mux/_018_ ;
wire \dpath/a_mux/_019_ ;
wire \dpath/a_mux/_020_ ;
wire \dpath/a_mux/_021_ ;
wire \dpath/a_mux/_022_ ;
wire \dpath/a_mux/_023_ ;
wire \dpath/a_mux/_024_ ;
wire \dpath/a_mux/_025_ ;
wire \dpath/a_mux/_026_ ;
wire \dpath/a_mux/_027_ ;
wire \dpath/a_mux/_028_ ;
wire \dpath/a_mux/_029_ ;
wire \dpath/a_mux/_030_ ;
wire \dpath/a_mux/_031_ ;
wire \dpath/a_mux/_032_ ;
wire \dpath/a_mux/_033_ ;
wire \dpath/a_mux/_034_ ;
wire \dpath/a_mux/_035_ ;
wire \dpath/a_mux/_036_ ;
wire \dpath/a_mux/_037_ ;
wire \dpath/a_mux/_038_ ;
wire \dpath/a_mux/_039_ ;
wire \dpath/a_mux/_040_ ;
wire \dpath/a_mux/_041_ ;
wire \dpath/a_mux/_042_ ;
wire \dpath/a_mux/_043_ ;
wire \dpath/a_mux/_044_ ;
wire \dpath/a_mux/_045_ ;
wire \dpath/a_mux/_046_ ;
wire \dpath/a_mux/_047_ ;
wire \dpath/a_mux/_048_ ;
wire \dpath/a_mux/_049_ ;
wire \dpath/a_mux/_050_ ;
wire \dpath/a_mux/_051_ ;
wire \dpath/a_mux/_052_ ;
wire \dpath/a_mux/_053_ ;
wire \dpath/a_mux/_054_ ;
wire \dpath/a_mux/_055_ ;
wire \dpath/a_mux/_056_ ;
wire \dpath/a_mux/_057_ ;
wire \dpath/a_mux/_058_ ;
wire \dpath/a_mux/_059_ ;
wire \dpath/a_mux/_060_ ;
wire \dpath/a_mux/_061_ ;
wire \dpath/a_mux/_062_ ;
wire \dpath/a_mux/_063_ ;
wire \dpath/a_mux/_064_ ;
wire \dpath/a_mux/_065_ ;
wire \dpath/a_mux/_066_ ;
wire \dpath/a_mux/_067_ ;
wire \dpath/a_mux/_068_ ;
wire \dpath/a_mux/_069_ ;
wire \dpath/a_mux/_070_ ;
wire \dpath/a_mux/_071_ ;
wire \dpath/a_mux/_072_ ;
wire \dpath/a_mux/_073_ ;
wire \dpath/a_mux/_074_ ;
wire \dpath/a_mux/_075_ ;
wire \dpath/a_mux/_076_ ;
wire \dpath/a_mux/_077_ ;
wire \dpath/a_mux/_078_ ;
wire \dpath/a_mux/_079_ ;
wire \dpath/a_mux/_080_ ;
wire \dpath/a_mux/_081_ ;
wire \dpath/a_mux/_082_ ;
wire \dpath/a_mux/_083_ ;
wire \dpath/a_mux/_084_ ;
wire \dpath/a_mux/_085_ ;
wire \dpath/a_mux/_086_ ;
wire \dpath/a_mux/_087_ ;
wire \dpath/a_mux/_088_ ;
wire \dpath/a_mux/_089_ ;
wire \dpath/a_mux/_090_ ;
wire \dpath/a_mux/_091_ ;
wire \dpath/a_mux/_092_ ;
wire \dpath/a_mux/_093_ ;
wire \dpath/a_mux/_094_ ;
wire \dpath/a_mux/_095_ ;
wire \dpath/a_mux/_096_ ;
wire \dpath/a_mux/_097_ ;
wire \dpath/a_mux/_098_ ;
wire \dpath/a_mux/_099_ ;
wire \dpath/a_mux/_100_ ;
wire \dpath/a_mux/_101_ ;
wire \dpath/a_mux/_102_ ;
wire \dpath/a_mux/_103_ ;
wire \dpath/a_mux/_104_ ;
wire \resp_msg[0] ;
wire \req_msg[16] ;
wire \resp_msg[1] ;
wire \req_msg[17] ;
wire \resp_msg[2] ;
wire \req_msg[18] ;
wire \resp_msg[3] ;
wire \req_msg[19] ;
wire \resp_msg[4] ;
wire \req_msg[20] ;
wire \resp_msg[5] ;
wire \req_msg[21] ;
wire \resp_msg[6] ;
wire \req_msg[22] ;
wire \resp_msg[7] ;
wire \req_msg[23] ;
wire \resp_msg[8] ;
wire \req_msg[24] ;
wire \resp_msg[9] ;
wire \req_msg[25] ;
wire \resp_msg[10] ;
wire \req_msg[26] ;
wire \resp_msg[11] ;
wire \req_msg[27] ;
wire \resp_msg[12] ;
wire \req_msg[28] ;
wire \resp_msg[13] ;
wire \req_msg[29] ;
wire \resp_msg[14] ;
wire \req_msg[30] ;
wire \resp_msg[15] ;
wire \req_msg[31] ;
wire \dpath/a_reg/_000_ ;
wire \dpath/a_reg/_001_ ;
wire \dpath/a_reg/_002_ ;
wire \dpath/a_reg/_003_ ;
wire \dpath/a_reg/_004_ ;
wire \dpath/a_reg/_005_ ;
wire \dpath/a_reg/_006_ ;
wire \dpath/a_reg/_007_ ;
wire \dpath/a_reg/_008_ ;
wire \dpath/a_reg/_009_ ;
wire \dpath/a_reg/_010_ ;
wire \dpath/a_reg/_011_ ;
wire \dpath/a_reg/_012_ ;
wire \dpath/a_reg/_013_ ;
wire \dpath/a_reg/_014_ ;
wire \dpath/a_reg/_015_ ;
wire \dpath/a_reg/_016_ ;
wire \dpath/a_reg/_017_ ;
wire \dpath/a_reg/_018_ ;
wire \dpath/a_reg/_019_ ;
wire \dpath/a_reg/_020_ ;
wire \dpath/a_reg/_021_ ;
wire \dpath/a_reg/_022_ ;
wire \dpath/a_reg/_023_ ;
wire \dpath/a_reg/_024_ ;
wire \dpath/a_reg/_025_ ;
wire \dpath/a_reg/_026_ ;
wire \dpath/a_reg/_027_ ;
wire \dpath/a_reg/_028_ ;
wire \dpath/a_reg/_029_ ;
wire \dpath/a_reg/_030_ ;
wire \dpath/a_reg/_031_ ;
wire \dpath/a_reg/_032_ ;
wire \dpath/a_reg/_033_ ;
wire \dpath/a_reg/_034_ ;
wire \dpath/a_reg/_035_ ;
wire \dpath/a_reg/_036_ ;
wire \dpath/a_reg/_037_ ;
wire \dpath/a_reg/_038_ ;
wire \dpath/a_reg/_039_ ;
wire \dpath/a_reg/_040_ ;
wire \dpath/a_reg/_041_ ;
wire \dpath/a_reg/_042_ ;
wire \dpath/a_reg/_043_ ;
wire \dpath/a_reg/_044_ ;
wire \dpath/a_reg/_045_ ;
wire \dpath/a_reg/_046_ ;
wire \dpath/a_reg/_047_ ;
wire \dpath/a_reg/_048_ ;
wire \dpath/a_reg/_049_ ;
wire \dpath/a_reg/_050_ ;
wire \dpath/a_reg/_051_ ;
wire \dpath/a_reg/_052_ ;
wire \dpath/a_reg/_053_ ;
wire \dpath/a_reg/_054_ ;
wire \dpath/a_reg/_055_ ;
wire \dpath/a_reg/_056_ ;
wire \dpath/a_reg/_057_ ;
wire \dpath/a_reg/_058_ ;
wire \dpath/a_reg/_059_ ;
wire \dpath/a_reg/_060_ ;
wire \dpath/a_reg/_061_ ;
wire \dpath/a_reg/_062_ ;
wire \dpath/a_reg/_063_ ;
wire \dpath/a_reg/_064_ ;
wire \dpath/a_reg/_065_ ;
wire \dpath/a_reg/_066_ ;
wire \dpath/a_reg/_067_ ;
wire \dpath/a_reg/_068_ ;
wire \dpath/a_reg/_069_ ;
wire \dpath/a_reg/_070_ ;
wire \dpath/a_reg/_071_ ;
wire \dpath/a_reg/_072_ ;
wire \dpath/a_reg/_073_ ;
wire \dpath/a_reg/_074_ ;
wire \dpath/a_reg/_075_ ;
wire \dpath/a_reg/_076_ ;
wire \dpath/a_reg/_077_ ;
wire \dpath/a_reg/_078_ ;
wire \dpath/a_reg/_079_ ;
wire \dpath/a_reg/_080_ ;
wire \dpath/b_mux/_000_ ;
wire \dpath/b_mux/_001_ ;
wire \dpath/b_mux/_002_ ;
wire \dpath/b_mux/_003_ ;
wire \dpath/b_mux/_004_ ;
wire \dpath/b_mux/_005_ ;
wire \dpath/b_mux/_006_ ;
wire \dpath/b_mux/_007_ ;
wire \dpath/b_mux/_008_ ;
wire \dpath/b_mux/_009_ ;
wire \dpath/b_mux/_010_ ;
wire \dpath/b_mux/_011_ ;
wire \dpath/b_mux/_012_ ;
wire \dpath/b_mux/_013_ ;
wire \dpath/b_mux/_014_ ;
wire \dpath/b_mux/_015_ ;
wire \dpath/b_mux/_016_ ;
wire \dpath/b_mux/_017_ ;
wire \dpath/b_mux/_018_ ;
wire \dpath/b_mux/_019_ ;
wire \dpath/b_mux/_020_ ;
wire \dpath/b_mux/_021_ ;
wire \dpath/b_mux/_022_ ;
wire \dpath/b_mux/_023_ ;
wire \dpath/b_mux/_024_ ;
wire \dpath/b_mux/_025_ ;
wire \dpath/b_mux/_026_ ;
wire \dpath/b_mux/_027_ ;
wire \dpath/b_mux/_028_ ;
wire \dpath/b_mux/_029_ ;
wire \dpath/b_mux/_030_ ;
wire \dpath/b_mux/_031_ ;
wire \dpath/b_mux/_032_ ;
wire \dpath/b_mux/_033_ ;
wire \dpath/b_mux/_034_ ;
wire \dpath/b_mux/_035_ ;
wire \dpath/b_mux/_036_ ;
wire \dpath/b_mux/_037_ ;
wire \dpath/b_mux/_038_ ;
wire \dpath/b_mux/_039_ ;
wire \dpath/b_mux/_040_ ;
wire \dpath/b_mux/_041_ ;
wire \dpath/b_mux/_042_ ;
wire \dpath/b_mux/_043_ ;
wire \dpath/b_mux/_044_ ;
wire \dpath/b_mux/_045_ ;
wire \dpath/b_mux/_046_ ;
wire \dpath/b_mux/_047_ ;
wire \dpath/b_mux/_048_ ;
wire \req_msg[0] ;
wire \req_msg[1] ;
wire \req_msg[2] ;
wire \req_msg[3] ;
wire \req_msg[4] ;
wire \req_msg[5] ;
wire \req_msg[6] ;
wire \req_msg[7] ;
wire \req_msg[8] ;
wire \req_msg[9] ;
wire \req_msg[10] ;
wire \req_msg[11] ;
wire \req_msg[12] ;
wire \req_msg[13] ;
wire \req_msg[14] ;
wire \req_msg[15] ;
wire \dpath/b_reg/_000_ ;
wire \dpath/b_reg/_001_ ;
wire \dpath/b_reg/_002_ ;
wire \dpath/b_reg/_003_ ;
wire \dpath/b_reg/_004_ ;
wire \dpath/b_reg/_005_ ;
wire \dpath/b_reg/_006_ ;
wire \dpath/b_reg/_007_ ;
wire \dpath/b_reg/_008_ ;
wire \dpath/b_reg/_009_ ;
wire \dpath/b_reg/_010_ ;
wire \dpath/b_reg/_011_ ;
wire \dpath/b_reg/_012_ ;
wire \dpath/b_reg/_013_ ;
wire \dpath/b_reg/_014_ ;
wire \dpath/b_reg/_015_ ;
wire \dpath/b_reg/_016_ ;
wire \dpath/b_reg/_017_ ;
wire \dpath/b_reg/_018_ ;
wire \dpath/b_reg/_019_ ;
wire \dpath/b_reg/_020_ ;
wire \dpath/b_reg/_021_ ;
wire \dpath/b_reg/_022_ ;
wire \dpath/b_reg/_023_ ;
wire \dpath/b_reg/_024_ ;
wire \dpath/b_reg/_025_ ;
wire \dpath/b_reg/_026_ ;
wire \dpath/b_reg/_027_ ;
wire \dpath/b_reg/_028_ ;
wire \dpath/b_reg/_029_ ;
wire \dpath/b_reg/_030_ ;
wire \dpath/b_reg/_031_ ;
wire \dpath/b_reg/_032_ ;
wire \dpath/b_reg/_033_ ;
wire \dpath/b_reg/_034_ ;
wire \dpath/b_reg/_035_ ;
wire \dpath/b_reg/_036_ ;
wire \dpath/b_reg/_037_ ;
wire \dpath/b_reg/_038_ ;
wire \dpath/b_reg/_039_ ;
wire \dpath/b_reg/_040_ ;
wire \dpath/b_reg/_041_ ;
wire \dpath/b_reg/_042_ ;
wire \dpath/b_reg/_043_ ;
wire \dpath/b_reg/_044_ ;
wire \dpath/b_reg/_045_ ;
wire \dpath/b_reg/_046_ ;
wire \dpath/b_reg/_047_ ;
wire \dpath/b_reg/_048_ ;
wire \dpath/b_reg/_049_ ;
wire \dpath/b_reg/_050_ ;
wire \dpath/b_reg/_051_ ;
wire \dpath/b_reg/_052_ ;
wire \dpath/b_reg/_053_ ;
wire \dpath/b_reg/_054_ ;
wire \dpath/b_reg/_055_ ;
wire \dpath/b_reg/_056_ ;
wire \dpath/b_reg/_057_ ;
wire \dpath/b_reg/_058_ ;
wire \dpath/b_reg/_059_ ;
wire \dpath/b_reg/_060_ ;
wire \dpath/b_reg/_061_ ;
wire \dpath/b_reg/_062_ ;
wire \dpath/b_reg/_063_ ;
wire \dpath/b_reg/_064_ ;
wire \dpath/b_reg/_065_ ;
wire \dpath/b_reg/_066_ ;
wire \dpath/b_reg/_067_ ;
wire \dpath/b_reg/_068_ ;
wire \dpath/b_reg/_069_ ;
wire \dpath/b_reg/_070_ ;
wire \dpath/b_reg/_071_ ;
wire \dpath/b_reg/_072_ ;
wire \dpath/b_reg/_073_ ;
wire \dpath/b_reg/_074_ ;
wire \dpath/b_reg/_075_ ;
wire \dpath/b_reg/_076_ ;
wire \dpath/b_reg/_077_ ;
wire \dpath/b_reg/_078_ ;
wire \dpath/b_reg/_079_ ;
wire \dpath/b_reg/_080_ ;
wire \dpath/b_zero/_00_ ;
wire \dpath/b_zero/_01_ ;
wire \dpath/b_zero/_02_ ;
wire \dpath/b_zero/_03_ ;
wire \dpath/b_zero/_04_ ;
wire \dpath/b_zero/_05_ ;
wire \dpath/b_zero/_06_ ;
wire \dpath/b_zero/_07_ ;
wire \dpath/b_zero/_08_ ;
wire \dpath/b_zero/_09_ ;
wire \dpath/b_zero/_10_ ;
wire \dpath/b_zero/_11_ ;
wire \dpath/b_zero/_12_ ;
wire \dpath/b_zero/_13_ ;
wire \dpath/b_zero/_14_ ;
wire \dpath/b_zero/_15_ ;
wire \dpath/b_zero/_16_ ;
wire \dpath/b_zero/_17_ ;
wire \dpath/b_zero/_18_ ;
wire \dpath/b_zero/_19_ ;
wire \dpath/b_zero/_20_ ;
wire \dpath/sub/_000_ ;
wire \dpath/sub/_001_ ;
wire \dpath/sub/_002_ ;
wire \dpath/sub/_003_ ;
wire \dpath/sub/_004_ ;
wire \dpath/sub/_005_ ;
wire \dpath/sub/_006_ ;
wire \dpath/sub/_007_ ;
wire \dpath/sub/_008_ ;
wire \dpath/sub/_009_ ;
wire \dpath/sub/_010_ ;
wire \dpath/sub/_011_ ;
wire \dpath/sub/_012_ ;
wire \dpath/sub/_013_ ;
wire \dpath/sub/_014_ ;
wire \dpath/sub/_015_ ;
wire \dpath/sub/_016_ ;
wire \dpath/sub/_017_ ;
wire \dpath/sub/_018_ ;
wire \dpath/sub/_019_ ;
wire \dpath/sub/_020_ ;
wire \dpath/sub/_021_ ;
wire \dpath/sub/_022_ ;
wire \dpath/sub/_023_ ;
wire \dpath/sub/_024_ ;
wire \dpath/sub/_025_ ;
wire \dpath/sub/_026_ ;
wire \dpath/sub/_027_ ;
wire \dpath/sub/_028_ ;
wire \dpath/sub/_029_ ;
wire \dpath/sub/_030_ ;
wire \dpath/sub/_031_ ;
wire \dpath/sub/_032_ ;
wire \dpath/sub/_033_ ;
wire \dpath/sub/_034_ ;
wire \dpath/sub/_035_ ;
wire \dpath/sub/_036_ ;
wire \dpath/sub/_037_ ;
wire \dpath/sub/_038_ ;
wire \dpath/sub/_039_ ;
wire \dpath/sub/_040_ ;
wire \dpath/sub/_041_ ;
wire \dpath/sub/_042_ ;
wire \dpath/sub/_043_ ;
wire \dpath/sub/_044_ ;
wire \dpath/sub/_045_ ;
wire \dpath/sub/_046_ ;
wire \dpath/sub/_047_ ;
wire \dpath/sub/_048_ ;
wire \dpath/sub/_049_ ;
wire \dpath/sub/_050_ ;
wire \dpath/sub/_051_ ;
wire \dpath/sub/_052_ ;
wire \dpath/sub/_053_ ;
wire \dpath/sub/_054_ ;
wire \dpath/sub/_055_ ;
wire \dpath/sub/_056_ ;
wire \dpath/sub/_057_ ;
wire \dpath/sub/_058_ ;
wire \dpath/sub/_059_ ;
wire \dpath/sub/_060_ ;
wire \dpath/sub/_061_ ;
wire \dpath/sub/_062_ ;
wire \dpath/sub/_063_ ;
wire \dpath/sub/_064_ ;
wire \dpath/sub/_065_ ;
wire \dpath/sub/_066_ ;
wire \dpath/sub/_067_ ;
wire \dpath/sub/_068_ ;
wire \dpath/sub/_069_ ;
wire \dpath/sub/_070_ ;
wire \dpath/sub/_071_ ;
wire \dpath/sub/_072_ ;
wire \dpath/sub/_073_ ;
wire \dpath/sub/_074_ ;
wire \dpath/sub/_075_ ;
wire \dpath/sub/_076_ ;
wire \dpath/sub/_077_ ;
wire \dpath/sub/_078_ ;
wire \dpath/sub/_079_ ;
wire \dpath/sub/_080_ ;
wire \dpath/sub/_081_ ;
wire \dpath/sub/_082_ ;
wire \dpath/sub/_083_ ;
wire \dpath/sub/_084_ ;
wire \dpath/sub/_085_ ;
wire \dpath/sub/_086_ ;
wire \dpath/sub/_087_ ;
wire \dpath/sub/_088_ ;
wire \dpath/sub/_089_ ;
wire \dpath/sub/_090_ ;
wire \dpath/sub/_091_ ;
wire \dpath/sub/_092_ ;
wire \dpath/sub/_093_ ;
wire \dpath/sub/_094_ ;
wire \dpath/sub/_095_ ;
wire \dpath/sub/_096_ ;
wire \dpath/sub/_097_ ;
wire \dpath/sub/_098_ ;
wire \dpath/sub/_099_ ;
wire \dpath/sub/_100_ ;
wire \dpath/sub/_101_ ;
wire \dpath/sub/_102_ ;
wire \dpath/sub/_103_ ;
wire \dpath/sub/_104_ ;
wire \dpath/sub/_105_ ;
wire \dpath/sub/_106_ ;
wire \dpath/sub/_107_ ;
wire \dpath/sub/_108_ ;
wire \dpath/sub/_109_ ;
wire \dpath/sub/_110_ ;
wire \dpath/sub/_111_ ;
wire \dpath/sub/_112_ ;
wire \dpath/sub/_113_ ;
wire \dpath/sub/_114_ ;
wire \dpath/sub/_115_ ;
wire \dpath/sub/_116_ ;
wire \dpath/sub/_117_ ;
wire \dpath/sub/_118_ ;
wire \dpath/sub/_119_ ;
wire \dpath/sub/_120_ ;
wire \dpath/sub/_121_ ;
wire \dpath/sub/_122_ ;
wire \dpath/sub/_123_ ;
wire \dpath/sub/_124_ ;
wire \dpath/sub/_125_ ;
wire \dpath/sub/_126_ ;
wire \dpath/sub/_127_ ;
wire \dpath/sub/_128_ ;
wire \dpath/sub/_129_ ;
wire \dpath/sub/_130_ ;
wire \dpath/sub/_131_ ;
wire \dpath/sub/_132_ ;
wire \dpath/sub/_133_ ;
wire \dpath/sub/_134_ ;
wire \dpath/sub/_135_ ;
wire \dpath/sub/_136_ ;
wire \dpath/sub/_137_ ;
wire \dpath/sub/_138_ ;
wire \dpath/sub/_139_ ;

NOR2_X1 \ctrl/_20_ ( .A1(\ctrl/_05_ ), .A2(\ctrl/_06_ ), .ZN(\ctrl/_03_ ) );
INV_X32 \ctrl/_21_ ( .A(\ctrl/_06_ ), .ZN(\ctrl/_02_ ) );
NOR2_X1 \ctrl/_22_ ( .A1(\ctrl/_02_ ), .A2(\ctrl/_05_ ), .ZN(\ctrl/_19_ ) );
INV_X32 \ctrl/_23_ ( .A(\ctrl/_05_ ), .ZN(\ctrl/_09_ ) );
NOR3_X1 \ctrl/_24_ ( .A1(\ctrl/_09_ ), .A2(\ctrl/_06_ ), .A3(\ctrl/_07_ ), .ZN(\ctrl/_00_ ) );
AND3_X4 \ctrl/_25_ ( .A1(\ctrl/_02_ ), .A2(\ctrl/_05_ ), .A3(\ctrl/_07_ ), .ZN(\ctrl/_01_ ) );
NOR2_X4 \ctrl/_26_ ( .A1(\ctrl/_09_ ), .A2(\ctrl/_06_ ), .ZN(\ctrl/_10_ ) );
INV_X8 \ctrl/_27_ ( .A(\ctrl/_07_ ), .ZN(\ctrl/_11_ ) );
AND3_X4 \ctrl/_28_ ( .A1(\ctrl/_10_ ), .A2(\ctrl/_11_ ), .A3(\ctrl/_08_ ), .ZN(\ctrl/_12_ ) );
NAND2_X1 \ctrl/_29_ ( .A1(\ctrl/_02_ ), .A2(\ctrl/_17_ ), .ZN(\ctrl/_13_ ) );
AOI21_X1 \ctrl/_30_ ( .A(\ctrl/_12_ ), .B1(\ctrl/_09_ ), .B2(\ctrl/_13_ ), .ZN(\ctrl/_15_ ) );
INV_X1 \ctrl/_31_ ( .A(\ctrl/_12_ ), .ZN(\ctrl/_14_ ) );
AOI22_X1 \ctrl/_32_ ( .A1(\ctrl/_14_ ), .A2(\ctrl/_02_ ), .B1(\ctrl/_18_ ), .B2(\ctrl/_19_ ), .ZN(\ctrl/_16_ ) );
AOI21_X1 \ctrl/_33_ ( .A(\ctrl/_06_ ), .B1(\ctrl/_11_ ), .B2(\ctrl/_05_ ), .ZN(\ctrl/_04_ ) );
BUF_X1 \ctrl/_34_ ( .A(ctrl$b_mux_sel ), .Z(req_rdy ) );
BUF_X1 \ctrl/_35_ ( .A(\ctrl/curr_state__0[0] ), .Z(\ctrl/_05_ ) );
BUF_X1 \ctrl/_36_ ( .A(\ctrl/curr_state__0[1] ), .Z(\ctrl/_06_ ) );
BUF_X1 \ctrl/_37_ ( .A(\ctrl/_03_ ), .Z(ctrl$b_mux_sel ) );
BUF_X1 \ctrl/_38_ ( .A(\ctrl/_19_ ), .Z(resp_val ) );
BUF_X1 \ctrl/_39_ ( .A(ctrl$is_a_lt_b ), .Z(\ctrl/_07_ ) );
BUF_X1 \ctrl/_40_ ( .A(\ctrl/_00_ ), .Z(\ctrl$a_mux_sel[0] ) );
BUF_X1 \ctrl/_41_ ( .A(\ctrl/_01_ ), .Z(\ctrl$a_mux_sel[1] ) );
BUF_X1 \ctrl/_42_ ( .A(req_val ), .Z(\ctrl/_17_ ) );
BUF_X1 \ctrl/_43_ ( .A(ctrl$is_b_zero ), .Z(\ctrl/_08_ ) );
BUF_X1 \ctrl/_44_ ( .A(resp_rdy ), .Z(\ctrl/_18_ ) );
BUF_X1 \ctrl/_45_ ( .A(\ctrl/_15_ ), .Z(\ctrl/next_state__0[0] ) );
BUF_X1 \ctrl/_46_ ( .A(\ctrl/_16_ ), .Z(\ctrl/next_state__0[1] ) );
BUF_X1 \ctrl/_47_ ( .A(\ctrl/_04_ ), .Z(ctrl$b_reg_en ) );
BUF_X1 \ctrl/_48_ ( .A(\ctrl/_02_ ), .Z(ctrl$a_reg_en ) );
INV_X16 \ctrl/state/_11_ ( .A(\ctrl/state/_04_ ), .ZN(\ctrl/state/_06_ ) );
NOR2_X1 \ctrl/state/_12_ ( .A1(\ctrl/state/_06_ ), .A2(\ctrl/state/_08_ ), .ZN(\ctrl/state/_02_ ) );
INV_X16 \ctrl/state/_13_ ( .A(\ctrl/state/_05_ ), .ZN(\ctrl/state/_07_ ) );
NOR2_X1 \ctrl/state/_14_ ( .A1(\ctrl/state/_07_ ), .A2(\ctrl/state/_08_ ), .ZN(\ctrl/state/_03_ ) );
BUF_X1 \ctrl/state/_15_ ( .A(\ctrl/next_state__0[0] ), .Z(\ctrl/state/_04_ ) );
BUF_X1 \ctrl/state/_16_ ( .A(reset ), .Z(\ctrl/state/_08_ ) );
BUF_X1 \ctrl/state/_17_ ( .A(\ctrl/state/_02_ ), .Z(\ctrl/state/_00_ ) );
BUF_X1 \ctrl/state/_18_ ( .A(\ctrl/next_state__0[1] ), .Z(\ctrl/state/_05_ ) );
BUF_X1 \ctrl/state/_19_ ( .A(\ctrl/state/_03_ ), .Z(\ctrl/state/_01_ ) );
DFF_X1 \ctrl/state/_20_ ( .CK(clk ), .D(\ctrl/state/_00_ ), .Q(\ctrl/curr_state__0[0] ), .QN(\ctrl/state/_09_ ) );
DFF_X1 \ctrl/state/_21_ ( .CK(clk ), .D(\ctrl/state/_01_ ), .Q(\ctrl/curr_state__0[1] ), .QN(\ctrl/state/_10_ ) );
XNOR2_X2 \dpath/a_lt_b/_109_ ( .A(\dpath/a_lt_b/_022_ ), .B(\dpath/a_lt_b/_006_ ), .ZN(\dpath/a_lt_b/_042_ ) );
INV_X2 \dpath/a_lt_b/_110_ ( .A(\dpath/a_lt_b/_042_ ), .ZN(\dpath/a_lt_b/_043_ ) );
INV_X16 \dpath/a_lt_b/_111_ ( .A(\dpath/a_lt_b/_021_ ), .ZN(\dpath/a_lt_b/_044_ ) );
NOR2_X1 \dpath/a_lt_b/_112_ ( .A1(\dpath/a_lt_b/_044_ ), .A2(\dpath/a_lt_b/_005_ ), .ZN(\dpath/a_lt_b/_045_ ) );
AND2_X2 \dpath/a_lt_b/_113_ ( .A1(\dpath/a_lt_b/_044_ ), .A2(\dpath/a_lt_b/_005_ ), .ZN(\dpath/a_lt_b/_046_ ) );
NOR3_X2 \dpath/a_lt_b/_114_ ( .A1(\dpath/a_lt_b/_043_ ), .A2(\dpath/a_lt_b/_045_ ), .A3(\dpath/a_lt_b/_046_ ), .ZN(\dpath/a_lt_b/_047_ ) );
INV_X1 \dpath/a_lt_b/_115_ ( .A(\dpath/a_lt_b/_003_ ), .ZN(\dpath/a_lt_b/_048_ ) );
NAND2_X1 \dpath/a_lt_b/_116_ ( .A1(\dpath/a_lt_b/_048_ ), .A2(\dpath/a_lt_b/_019_ ), .ZN(\dpath/a_lt_b/_049_ ) );
INV_X1 \dpath/a_lt_b/_117_ ( .A(\dpath/a_lt_b/_020_ ), .ZN(\dpath/a_lt_b/_050_ ) );
OAI21_X1 \dpath/a_lt_b/_118_ ( .A(\dpath/a_lt_b/_049_ ), .B1(\dpath/a_lt_b/_004_ ), .B2(\dpath/a_lt_b/_050_ ), .ZN(\dpath/a_lt_b/_051_ ) );
NAND2_X1 \dpath/a_lt_b/_119_ ( .A1(\dpath/a_lt_b/_050_ ), .A2(\dpath/a_lt_b/_004_ ), .ZN(\dpath/a_lt_b/_052_ ) );
OAI21_X1 \dpath/a_lt_b/_120_ ( .A(\dpath/a_lt_b/_052_ ), .B1(\dpath/a_lt_b/_019_ ), .B2(\dpath/a_lt_b/_048_ ), .ZN(\dpath/a_lt_b/_053_ ) );
NOR2_X1 \dpath/a_lt_b/_121_ ( .A1(\dpath/a_lt_b/_051_ ), .A2(\dpath/a_lt_b/_053_ ), .ZN(\dpath/a_lt_b/_054_ ) );
AND2_X2 \dpath/a_lt_b/_122_ ( .A1(\dpath/a_lt_b/_047_ ), .A2(\dpath/a_lt_b/_054_ ), .ZN(\dpath/a_lt_b/_055_ ) );
INV_X32 \dpath/a_lt_b/_123_ ( .A(\dpath/a_lt_b/_018_ ), .ZN(\dpath/a_lt_b/_056_ ) );
NOR2_X4 \dpath/a_lt_b/_124_ ( .A1(\dpath/a_lt_b/_056_ ), .A2(\dpath/a_lt_b/_002_ ), .ZN(\dpath/a_lt_b/_057_ ) );
INV_X32 \dpath/a_lt_b/_125_ ( .A(\dpath/a_lt_b/_017_ ), .ZN(\dpath/a_lt_b/_058_ ) );
AOI21_X1 \dpath/a_lt_b/_126_ ( .A(\dpath/a_lt_b/_057_ ), .B1(\dpath/a_lt_b/_058_ ), .B2(\dpath/a_lt_b/_001_ ), .ZN(\dpath/a_lt_b/_059_ ) );
NOR2_X4 \dpath/a_lt_b/_127_ ( .A1(\dpath/a_lt_b/_058_ ), .A2(\dpath/a_lt_b/_001_ ), .ZN(\dpath/a_lt_b/_060_ ) );
AOI21_X1 \dpath/a_lt_b/_128_ ( .A(\dpath/a_lt_b/_060_ ), .B1(\dpath/a_lt_b/_002_ ), .B2(\dpath/a_lt_b/_056_ ), .ZN(\dpath/a_lt_b/_061_ ) );
AND2_X2 \dpath/a_lt_b/_129_ ( .A1(\dpath/a_lt_b/_059_ ), .A2(\dpath/a_lt_b/_061_ ), .ZN(\dpath/a_lt_b/_062_ ) );
XOR2_X1 \dpath/a_lt_b/_130_ ( .A(\dpath/a_lt_b/_030_ ), .B(\dpath/a_lt_b/_014_ ), .Z(\dpath/a_lt_b/_063_ ) );
INV_X32 \dpath/a_lt_b/_131_ ( .A(\dpath/a_lt_b/_031_ ), .ZN(\dpath/a_lt_b/_064_ ) );
NOR2_X1 \dpath/a_lt_b/_132_ ( .A1(\dpath/a_lt_b/_064_ ), .A2(\dpath/a_lt_b/_015_ ), .ZN(\dpath/a_lt_b/_065_ ) );
AND2_X1 \dpath/a_lt_b/_133_ ( .A1(\dpath/a_lt_b/_064_ ), .A2(\dpath/a_lt_b/_015_ ), .ZN(\dpath/a_lt_b/_066_ ) );
NOR3_X1 \dpath/a_lt_b/_134_ ( .A1(\dpath/a_lt_b/_063_ ), .A2(\dpath/a_lt_b/_065_ ), .A3(\dpath/a_lt_b/_066_ ), .ZN(\dpath/a_lt_b/_067_ ) );
AND3_X2 \dpath/a_lt_b/_135_ ( .A1(\dpath/a_lt_b/_055_ ), .A2(\dpath/a_lt_b/_062_ ), .A3(\dpath/a_lt_b/_067_ ), .ZN(\dpath/a_lt_b/_068_ ) );
XOR2_X1 \dpath/a_lt_b/_136_ ( .A(\dpath/a_lt_b/_023_ ), .B(\dpath/a_lt_b/_007_ ), .Z(\dpath/a_lt_b/_069_ ) );
INV_X1 \dpath/a_lt_b/_137_ ( .A(\dpath/a_lt_b/_016_ ), .ZN(\dpath/a_lt_b/_070_ ) );
AOI21_X1 \dpath/a_lt_b/_138_ ( .A(\dpath/a_lt_b/_069_ ), .B1(\dpath/a_lt_b/_070_ ), .B2(\dpath/a_lt_b/_000_ ), .ZN(\dpath/a_lt_b/_071_ ) );
OAI211_X2 \dpath/a_lt_b/_139_ ( .A(\dpath/a_lt_b/_068_ ), .B(\dpath/a_lt_b/_071_ ), .C1(\dpath/a_lt_b/_070_ ), .C2(\dpath/a_lt_b/_000_ ), .ZN(\dpath/a_lt_b/_072_ ) );
INV_X2 \dpath/a_lt_b/_140_ ( .A(\dpath/a_lt_b/_013_ ), .ZN(\dpath/a_lt_b/_073_ ) );
OR2_X4 \dpath/a_lt_b/_141_ ( .A1(\dpath/a_lt_b/_073_ ), .A2(\dpath/a_lt_b/_029_ ), .ZN(\dpath/a_lt_b/_074_ ) );
NAND2_X1 \dpath/a_lt_b/_142_ ( .A1(\dpath/a_lt_b/_073_ ), .A2(\dpath/a_lt_b/_029_ ), .ZN(\dpath/a_lt_b/_075_ ) );
INV_X2 \dpath/a_lt_b/_143_ ( .A(\dpath/a_lt_b/_012_ ), .ZN(\dpath/a_lt_b/_076_ ) );
OAI211_X2 \dpath/a_lt_b/_144_ ( .A(\dpath/a_lt_b/_074_ ), .B(\dpath/a_lt_b/_075_ ), .C1(\dpath/a_lt_b/_028_ ), .C2(\dpath/a_lt_b/_076_ ), .ZN(\dpath/a_lt_b/_077_ ) );
AOI21_X2 \dpath/a_lt_b/_145_ ( .A(\dpath/a_lt_b/_077_ ), .B1(\dpath/a_lt_b/_028_ ), .B2(\dpath/a_lt_b/_076_ ), .ZN(\dpath/a_lt_b/_078_ ) );
INV_X1 \dpath/a_lt_b/_146_ ( .A(\dpath/a_lt_b/_011_ ), .ZN(\dpath/a_lt_b/_079_ ) );
AND2_X1 \dpath/a_lt_b/_147_ ( .A1(\dpath/a_lt_b/_079_ ), .A2(\dpath/a_lt_b/_027_ ), .ZN(\dpath/a_lt_b/_080_ ) );
INV_X1 \dpath/a_lt_b/_148_ ( .A(\dpath/a_lt_b/_010_ ), .ZN(\dpath/a_lt_b/_081_ ) );
AND2_X1 \dpath/a_lt_b/_149_ ( .A1(\dpath/a_lt_b/_081_ ), .A2(\dpath/a_lt_b/_026_ ), .ZN(\dpath/a_lt_b/_082_ ) );
NOR2_X1 \dpath/a_lt_b/_150_ ( .A1(\dpath/a_lt_b/_079_ ), .A2(\dpath/a_lt_b/_027_ ), .ZN(\dpath/a_lt_b/_083_ ) );
NOR2_X1 \dpath/a_lt_b/_151_ ( .A1(\dpath/a_lt_b/_081_ ), .A2(\dpath/a_lt_b/_026_ ), .ZN(\dpath/a_lt_b/_084_ ) );
NOR4_X4 \dpath/a_lt_b/_152_ ( .A1(\dpath/a_lt_b/_080_ ), .A2(\dpath/a_lt_b/_082_ ), .A3(\dpath/a_lt_b/_083_ ), .A4(\dpath/a_lt_b/_084_ ), .ZN(\dpath/a_lt_b/_085_ ) );
XNOR2_X1 \dpath/a_lt_b/_153_ ( .A(\dpath/a_lt_b/_025_ ), .B(\dpath/a_lt_b/_009_ ), .ZN(\dpath/a_lt_b/_086_ ) );
XNOR2_X1 \dpath/a_lt_b/_154_ ( .A(\dpath/a_lt_b/_024_ ), .B(\dpath/a_lt_b/_008_ ), .ZN(\dpath/a_lt_b/_087_ ) );
AND2_X1 \dpath/a_lt_b/_155_ ( .A1(\dpath/a_lt_b/_086_ ), .A2(\dpath/a_lt_b/_087_ ), .ZN(\dpath/a_lt_b/_088_ ) );
NAND3_X1 \dpath/a_lt_b/_156_ ( .A1(\dpath/a_lt_b/_078_ ), .A2(\dpath/a_lt_b/_085_ ), .A3(\dpath/a_lt_b/_088_ ), .ZN(\dpath/a_lt_b/_089_ ) );
NOR2_X2 \dpath/a_lt_b/_157_ ( .A1(\dpath/a_lt_b/_072_ ), .A2(\dpath/a_lt_b/_089_ ), .ZN(\dpath/a_lt_b/_090_ ) );
INV_X2 \dpath/a_lt_b/_158_ ( .A(\dpath/a_lt_b/_062_ ), .ZN(\dpath/a_lt_b/_091_ ) );
INV_X1 \dpath/a_lt_b/_159_ ( .A(\dpath/a_lt_b/_014_ ), .ZN(\dpath/a_lt_b/_092_ ) );
AOI21_X4 \dpath/a_lt_b/_160_ ( .A(\dpath/a_lt_b/_065_ ), .B1(\dpath/a_lt_b/_030_ ), .B2(\dpath/a_lt_b/_092_ ), .ZN(\dpath/a_lt_b/_093_ ) );
NOR3_X2 \dpath/a_lt_b/_161_ ( .A1(\dpath/a_lt_b/_091_ ), .A2(\dpath/a_lt_b/_093_ ), .A3(\dpath/a_lt_b/_066_ ), .ZN(\dpath/a_lt_b/_094_ ) );
AOI211_X4 \dpath/a_lt_b/_162_ ( .A(\dpath/a_lt_b/_001_ ), .B(\dpath/a_lt_b/_058_ ), .C1(\dpath/a_lt_b/_002_ ), .C2(\dpath/a_lt_b/_056_ ), .ZN(\dpath/a_lt_b/_095_ ) );
OR3_X2 \dpath/a_lt_b/_163_ ( .A1(\dpath/a_lt_b/_094_ ), .A2(\dpath/a_lt_b/_057_ ), .A3(\dpath/a_lt_b/_095_ ), .ZN(\dpath/a_lt_b/_096_ ) );
AND2_X2 \dpath/a_lt_b/_164_ ( .A1(\dpath/a_lt_b/_096_ ), .A2(\dpath/a_lt_b/_055_ ), .ZN(\dpath/a_lt_b/_097_ ) );
INV_X1 \dpath/a_lt_b/_165_ ( .A(\dpath/a_lt_b/_022_ ), .ZN(\dpath/a_lt_b/_098_ ) );
NOR2_X1 \dpath/a_lt_b/_166_ ( .A1(\dpath/a_lt_b/_098_ ), .A2(\dpath/a_lt_b/_006_ ), .ZN(\dpath/a_lt_b/_099_ ) );
AND3_X1 \dpath/a_lt_b/_167_ ( .A1(\dpath/a_lt_b/_047_ ), .A2(\dpath/a_lt_b/_051_ ), .A3(\dpath/a_lt_b/_052_ ), .ZN(\dpath/a_lt_b/_100_ ) );
AND2_X1 \dpath/a_lt_b/_168_ ( .A1(\dpath/a_lt_b/_042_ ), .A2(\dpath/a_lt_b/_045_ ), .ZN(\dpath/a_lt_b/_101_ ) );
NOR4_X4 \dpath/a_lt_b/_169_ ( .A1(\dpath/a_lt_b/_097_ ), .A2(\dpath/a_lt_b/_099_ ), .A3(\dpath/a_lt_b/_100_ ), .A4(\dpath/a_lt_b/_101_ ), .ZN(\dpath/a_lt_b/_102_ ) );
AOI211_X2 \dpath/a_lt_b/_170_ ( .A(\dpath/a_lt_b/_083_ ), .B(\dpath/a_lt_b/_077_ ), .C1(\dpath/a_lt_b/_028_ ), .C2(\dpath/a_lt_b/_076_ ), .ZN(\dpath/a_lt_b/_103_ ) );
OAI21_X1 \dpath/a_lt_b/_171_ ( .A(\dpath/a_lt_b/_103_ ), .B1(\dpath/a_lt_b/_080_ ), .B2(\dpath/a_lt_b/_082_ ), .ZN(\dpath/a_lt_b/_104_ ) );
NAND4_X1 \dpath/a_lt_b/_172_ ( .A1(\dpath/a_lt_b/_074_ ), .A2(\dpath/a_lt_b/_028_ ), .A3(\dpath/a_lt_b/_076_ ), .A4(\dpath/a_lt_b/_075_ ), .ZN(\dpath/a_lt_b/_105_ ) );
NAND3_X1 \dpath/a_lt_b/_173_ ( .A1(\dpath/a_lt_b/_104_ ), .A2(\dpath/a_lt_b/_075_ ), .A3(\dpath/a_lt_b/_105_ ), .ZN(\dpath/a_lt_b/_106_ ) );
NAND2_X1 \dpath/a_lt_b/_174_ ( .A1(\dpath/a_lt_b/_078_ ), .A2(\dpath/a_lt_b/_085_ ), .ZN(\dpath/a_lt_b/_107_ ) );
INV_X1 \dpath/a_lt_b/_175_ ( .A(\dpath/a_lt_b/_007_ ), .ZN(\dpath/a_lt_b/_032_ ) );
AND2_X1 \dpath/a_lt_b/_176_ ( .A1(\dpath/a_lt_b/_032_ ), .A2(\dpath/a_lt_b/_023_ ), .ZN(\dpath/a_lt_b/_033_ ) );
OAI21_X1 \dpath/a_lt_b/_177_ ( .A(\dpath/a_lt_b/_088_ ), .B1(\dpath/a_lt_b/_071_ ), .B2(\dpath/a_lt_b/_033_ ), .ZN(\dpath/a_lt_b/_034_ ) );
INV_X1 \dpath/a_lt_b/_178_ ( .A(\dpath/a_lt_b/_024_ ), .ZN(\dpath/a_lt_b/_035_ ) );
NOR2_X1 \dpath/a_lt_b/_179_ ( .A1(\dpath/a_lt_b/_035_ ), .A2(\dpath/a_lt_b/_008_ ), .ZN(\dpath/a_lt_b/_036_ ) );
AND2_X1 \dpath/a_lt_b/_180_ ( .A1(\dpath/a_lt_b/_086_ ), .A2(\dpath/a_lt_b/_036_ ), .ZN(\dpath/a_lt_b/_037_ ) );
INV_X1 \dpath/a_lt_b/_181_ ( .A(\dpath/a_lt_b/_009_ ), .ZN(\dpath/a_lt_b/_038_ ) );
AOI21_X1 \dpath/a_lt_b/_182_ ( .A(\dpath/a_lt_b/_037_ ), .B1(\dpath/a_lt_b/_025_ ), .B2(\dpath/a_lt_b/_038_ ), .ZN(\dpath/a_lt_b/_039_ ) );
AOI21_X2 \dpath/a_lt_b/_183_ ( .A(\dpath/a_lt_b/_107_ ), .B1(\dpath/a_lt_b/_034_ ), .B2(\dpath/a_lt_b/_039_ ), .ZN(\dpath/a_lt_b/_040_ ) );
OAI21_X1 \dpath/a_lt_b/_184_ ( .A(\dpath/a_lt_b/_068_ ), .B1(\dpath/a_lt_b/_106_ ), .B2(\dpath/a_lt_b/_040_ ), .ZN(\dpath/a_lt_b/_041_ ) );
AOI21_X1 \dpath/a_lt_b/_185_ ( .A(\dpath/a_lt_b/_090_ ), .B1(\dpath/a_lt_b/_102_ ), .B2(\dpath/a_lt_b/_041_ ), .ZN(\dpath/a_lt_b/_108_ ) );
BUF_X1 \dpath/a_lt_b/_186_ ( .A(\dpath/a_lt_b$in1[14] ), .Z(\dpath/a_lt_b/_021_ ) );
BUF_X1 \dpath/a_lt_b/_187_ ( .A(\dpath/a_lt_b$in0[14] ), .Z(\dpath/a_lt_b/_005_ ) );
BUF_X1 \dpath/a_lt_b/_188_ ( .A(\dpath/a_lt_b$in0[13] ), .Z(\dpath/a_lt_b/_004_ ) );
BUF_X1 \dpath/a_lt_b/_189_ ( .A(\dpath/a_lt_b$in1[13] ), .Z(\dpath/a_lt_b/_020_ ) );
BUF_X1 \dpath/a_lt_b/_190_ ( .A(\dpath/a_lt_b$in1[12] ), .Z(\dpath/a_lt_b/_019_ ) );
BUF_X1 \dpath/a_lt_b/_191_ ( .A(\dpath/a_lt_b$in0[12] ), .Z(\dpath/a_lt_b/_003_ ) );
BUF_X1 \dpath/a_lt_b/_192_ ( .A(\dpath/a_lt_b$in0[11] ), .Z(\dpath/a_lt_b/_002_ ) );
BUF_X1 \dpath/a_lt_b/_193_ ( .A(\dpath/a_lt_b$in1[11] ), .Z(\dpath/a_lt_b/_018_ ) );
BUF_X1 \dpath/a_lt_b/_194_ ( .A(\dpath/a_lt_b$in1[10] ), .Z(\dpath/a_lt_b/_017_ ) );
BUF_X1 \dpath/a_lt_b/_195_ ( .A(\dpath/a_lt_b$in0[10] ), .Z(\dpath/a_lt_b/_001_ ) );
BUF_X1 \dpath/a_lt_b/_196_ ( .A(\dpath/a_lt_b$in0[9] ), .Z(\dpath/a_lt_b/_015_ ) );
BUF_X1 \dpath/a_lt_b/_197_ ( .A(\dpath/a_lt_b$in1[9] ), .Z(\dpath/a_lt_b/_031_ ) );
BUF_X1 \dpath/a_lt_b/_198_ ( .A(\dpath/a_lt_b$in1[8] ), .Z(\dpath/a_lt_b/_030_ ) );
BUF_X1 \dpath/a_lt_b/_199_ ( .A(\dpath/a_lt_b$in0[8] ), .Z(\dpath/a_lt_b/_014_ ) );
BUF_X1 \dpath/a_lt_b/_200_ ( .A(\dpath/a_lt_b$in1[7] ), .Z(\dpath/a_lt_b/_029_ ) );
BUF_X1 \dpath/a_lt_b/_201_ ( .A(\dpath/a_lt_b$in0[7] ), .Z(\dpath/a_lt_b/_013_ ) );
BUF_X1 \dpath/a_lt_b/_202_ ( .A(\dpath/a_lt_b$in1[6] ), .Z(\dpath/a_lt_b/_028_ ) );
BUF_X1 \dpath/a_lt_b/_203_ ( .A(\dpath/a_lt_b$in0[6] ), .Z(\dpath/a_lt_b/_012_ ) );
BUF_X1 \dpath/a_lt_b/_204_ ( .A(\dpath/a_lt_b$in0[5] ), .Z(\dpath/a_lt_b/_011_ ) );
BUF_X1 \dpath/a_lt_b/_205_ ( .A(\dpath/a_lt_b$in1[5] ), .Z(\dpath/a_lt_b/_027_ ) );
BUF_X1 \dpath/a_lt_b/_206_ ( .A(\dpath/a_lt_b$in1[4] ), .Z(\dpath/a_lt_b/_026_ ) );
BUF_X1 \dpath/a_lt_b/_207_ ( .A(\dpath/a_lt_b$in0[4] ), .Z(\dpath/a_lt_b/_010_ ) );
BUF_X1 \dpath/a_lt_b/_208_ ( .A(\dpath/a_lt_b$in1[3] ), .Z(\dpath/a_lt_b/_025_ ) );
BUF_X1 \dpath/a_lt_b/_209_ ( .A(\dpath/a_lt_b$in0[3] ), .Z(\dpath/a_lt_b/_009_ ) );
BUF_X1 \dpath/a_lt_b/_210_ ( .A(\dpath/a_lt_b$in1[2] ), .Z(\dpath/a_lt_b/_024_ ) );
BUF_X1 \dpath/a_lt_b/_211_ ( .A(\dpath/a_lt_b$in0[2] ), .Z(\dpath/a_lt_b/_008_ ) );
BUF_X1 \dpath/a_lt_b/_212_ ( .A(\dpath/a_lt_b$in1[1] ), .Z(\dpath/a_lt_b/_023_ ) );
BUF_X1 \dpath/a_lt_b/_213_ ( .A(\dpath/a_lt_b$in0[1] ), .Z(\dpath/a_lt_b/_007_ ) );
BUF_X1 \dpath/a_lt_b/_214_ ( .A(\dpath/a_lt_b$in1[0] ), .Z(\dpath/a_lt_b/_016_ ) );
BUF_X1 \dpath/a_lt_b/_215_ ( .A(\dpath/a_lt_b$in0[0] ), .Z(\dpath/a_lt_b/_000_ ) );
BUF_X1 \dpath/a_lt_b/_216_ ( .A(\dpath/a_lt_b/_108_ ), .Z(ctrl$is_a_lt_b ) );
BUF_X1 \dpath/a_lt_b/_217_ ( .A(\dpath/a_lt_b$in1[15] ), .Z(\dpath/a_lt_b/_022_ ) );
BUF_X1 \dpath/a_lt_b/_218_ ( .A(\dpath/a_lt_b$in0[15] ), .Z(\dpath/a_lt_b/_006_ ) );
INV_X32 \dpath/a_mux/_105_ ( .A(\dpath/a_mux/_104_ ), .ZN(\dpath/a_mux/_062_ ) );
AND2_X2 \dpath/a_mux/_106_ ( .A1(\dpath/a_mux/_062_ ), .A2(\dpath/a_mux/_103_ ), .ZN(\dpath/a_mux/_063_ ) );
BUF_X8 \dpath/a_mux/_107_ ( .A(\dpath/a_mux/_063_ ), .Z(\dpath/a_mux/_064_ ) );
NOR2_X4 \dpath/a_mux/_108_ ( .A1(\dpath/a_mux/_062_ ), .A2(\dpath/a_mux/_103_ ), .ZN(\dpath/a_mux/_065_ ) );
BUF_X4 \dpath/a_mux/_109_ ( .A(\dpath/a_mux/_065_ ), .Z(\dpath/a_mux/_066_ ) );
AOI22_X1 \dpath/a_mux/_110_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_016_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_032_ ), .ZN(\dpath/a_mux/_067_ ) );
XNOR2_X2 \dpath/a_mux/_111_ ( .A(\dpath/a_mux/_103_ ), .B(\dpath/a_mux/_104_ ), .ZN(\dpath/a_mux/_068_ ) );
BUF_X4 \dpath/a_mux/_112_ ( .A(\dpath/a_mux/_068_ ), .Z(\dpath/a_mux/_069_ ) );
NAND2_X1 \dpath/a_mux/_113_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_000_ ), .ZN(\dpath/a_mux/_070_ ) );
NAND2_X1 \dpath/a_mux/_114_ ( .A1(\dpath/a_mux/_067_ ), .A2(\dpath/a_mux/_070_ ), .ZN(\dpath/a_mux/_087_ ) );
AOI22_X1 \dpath/a_mux/_115_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_023_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_039_ ), .ZN(\dpath/a_mux/_071_ ) );
NAND2_X1 \dpath/a_mux/_116_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_007_ ), .ZN(\dpath/a_mux/_072_ ) );
NAND2_X1 \dpath/a_mux/_117_ ( .A1(\dpath/a_mux/_071_ ), .A2(\dpath/a_mux/_072_ ), .ZN(\dpath/a_mux/_094_ ) );
AOI22_X1 \dpath/a_mux/_118_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_024_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_040_ ), .ZN(\dpath/a_mux/_073_ ) );
NAND2_X1 \dpath/a_mux/_119_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_008_ ), .ZN(\dpath/a_mux/_074_ ) );
NAND2_X1 \dpath/a_mux/_120_ ( .A1(\dpath/a_mux/_073_ ), .A2(\dpath/a_mux/_074_ ), .ZN(\dpath/a_mux/_095_ ) );
AOI22_X1 \dpath/a_mux/_121_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_025_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_041_ ), .ZN(\dpath/a_mux/_075_ ) );
NAND2_X1 \dpath/a_mux/_122_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_009_ ), .ZN(\dpath/a_mux/_076_ ) );
NAND2_X1 \dpath/a_mux/_123_ ( .A1(\dpath/a_mux/_075_ ), .A2(\dpath/a_mux/_076_ ), .ZN(\dpath/a_mux/_096_ ) );
AOI22_X1 \dpath/a_mux/_124_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_026_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_042_ ), .ZN(\dpath/a_mux/_077_ ) );
NAND2_X1 \dpath/a_mux/_125_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_010_ ), .ZN(\dpath/a_mux/_078_ ) );
NAND2_X1 \dpath/a_mux/_126_ ( .A1(\dpath/a_mux/_077_ ), .A2(\dpath/a_mux/_078_ ), .ZN(\dpath/a_mux/_097_ ) );
AOI22_X1 \dpath/a_mux/_127_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_027_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_043_ ), .ZN(\dpath/a_mux/_079_ ) );
NAND2_X1 \dpath/a_mux/_128_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_011_ ), .ZN(\dpath/a_mux/_080_ ) );
NAND2_X1 \dpath/a_mux/_129_ ( .A1(\dpath/a_mux/_079_ ), .A2(\dpath/a_mux/_080_ ), .ZN(\dpath/a_mux/_098_ ) );
AOI22_X1 \dpath/a_mux/_130_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_028_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_044_ ), .ZN(\dpath/a_mux/_081_ ) );
NAND2_X1 \dpath/a_mux/_131_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_012_ ), .ZN(\dpath/a_mux/_082_ ) );
NAND2_X1 \dpath/a_mux/_132_ ( .A1(\dpath/a_mux/_081_ ), .A2(\dpath/a_mux/_082_ ), .ZN(\dpath/a_mux/_099_ ) );
AOI22_X1 \dpath/a_mux/_133_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_029_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_045_ ), .ZN(\dpath/a_mux/_083_ ) );
NAND2_X1 \dpath/a_mux/_134_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_013_ ), .ZN(\dpath/a_mux/_084_ ) );
NAND2_X1 \dpath/a_mux/_135_ ( .A1(\dpath/a_mux/_083_ ), .A2(\dpath/a_mux/_084_ ), .ZN(\dpath/a_mux/_100_ ) );
AOI22_X1 \dpath/a_mux/_136_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_030_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_046_ ), .ZN(\dpath/a_mux/_085_ ) );
NAND2_X1 \dpath/a_mux/_137_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_014_ ), .ZN(\dpath/a_mux/_086_ ) );
NAND2_X1 \dpath/a_mux/_138_ ( .A1(\dpath/a_mux/_085_ ), .A2(\dpath/a_mux/_086_ ), .ZN(\dpath/a_mux/_101_ ) );
AOI22_X1 \dpath/a_mux/_139_ ( .A1(\dpath/a_mux/_064_ ), .A2(\dpath/a_mux/_031_ ), .B1(\dpath/a_mux/_066_ ), .B2(\dpath/a_mux/_047_ ), .ZN(\dpath/a_mux/_048_ ) );
NAND2_X2 \dpath/a_mux/_140_ ( .A1(\dpath/a_mux/_069_ ), .A2(\dpath/a_mux/_015_ ), .ZN(\dpath/a_mux/_049_ ) );
NAND2_X1 \dpath/a_mux/_141_ ( .A1(\dpath/a_mux/_048_ ), .A2(\dpath/a_mux/_049_ ), .ZN(\dpath/a_mux/_102_ ) );
AOI22_X1 \dpath/a_mux/_142_ ( .A1(\dpath/a_mux/_063_ ), .A2(\dpath/a_mux/_017_ ), .B1(\dpath/a_mux/_065_ ), .B2(\dpath/a_mux/_033_ ), .ZN(\dpath/a_mux/_050_ ) );
NAND2_X1 \dpath/a_mux/_143_ ( .A1(\dpath/a_mux/_068_ ), .A2(\dpath/a_mux/_001_ ), .ZN(\dpath/a_mux/_051_ ) );
NAND2_X1 \dpath/a_mux/_144_ ( .A1(\dpath/a_mux/_050_ ), .A2(\dpath/a_mux/_051_ ), .ZN(\dpath/a_mux/_088_ ) );
AOI22_X1 \dpath/a_mux/_145_ ( .A1(\dpath/a_mux/_063_ ), .A2(\dpath/a_mux/_018_ ), .B1(\dpath/a_mux/_065_ ), .B2(\dpath/a_mux/_034_ ), .ZN(\dpath/a_mux/_052_ ) );
NAND2_X1 \dpath/a_mux/_146_ ( .A1(\dpath/a_mux/_068_ ), .A2(\dpath/a_mux/_002_ ), .ZN(\dpath/a_mux/_053_ ) );
NAND2_X1 \dpath/a_mux/_147_ ( .A1(\dpath/a_mux/_052_ ), .A2(\dpath/a_mux/_053_ ), .ZN(\dpath/a_mux/_089_ ) );
AOI22_X1 \dpath/a_mux/_148_ ( .A1(\dpath/a_mux/_063_ ), .A2(\dpath/a_mux/_019_ ), .B1(\dpath/a_mux/_065_ ), .B2(\dpath/a_mux/_035_ ), .ZN(\dpath/a_mux/_054_ ) );
NAND2_X1 \dpath/a_mux/_149_ ( .A1(\dpath/a_mux/_068_ ), .A2(\dpath/a_mux/_003_ ), .ZN(\dpath/a_mux/_055_ ) );
NAND2_X1 \dpath/a_mux/_150_ ( .A1(\dpath/a_mux/_054_ ), .A2(\dpath/a_mux/_055_ ), .ZN(\dpath/a_mux/_090_ ) );
AOI22_X1 \dpath/a_mux/_151_ ( .A1(\dpath/a_mux/_063_ ), .A2(\dpath/a_mux/_020_ ), .B1(\dpath/a_mux/_065_ ), .B2(\dpath/a_mux/_036_ ), .ZN(\dpath/a_mux/_056_ ) );
NAND2_X1 \dpath/a_mux/_152_ ( .A1(\dpath/a_mux/_068_ ), .A2(\dpath/a_mux/_004_ ), .ZN(\dpath/a_mux/_057_ ) );
NAND2_X1 \dpath/a_mux/_153_ ( .A1(\dpath/a_mux/_056_ ), .A2(\dpath/a_mux/_057_ ), .ZN(\dpath/a_mux/_091_ ) );
AOI22_X1 \dpath/a_mux/_154_ ( .A1(\dpath/a_mux/_063_ ), .A2(\dpath/a_mux/_021_ ), .B1(\dpath/a_mux/_065_ ), .B2(\dpath/a_mux/_037_ ), .ZN(\dpath/a_mux/_058_ ) );
NAND2_X1 \dpath/a_mux/_155_ ( .A1(\dpath/a_mux/_068_ ), .A2(\dpath/a_mux/_005_ ), .ZN(\dpath/a_mux/_059_ ) );
NAND2_X1 \dpath/a_mux/_156_ ( .A1(\dpath/a_mux/_058_ ), .A2(\dpath/a_mux/_059_ ), .ZN(\dpath/a_mux/_092_ ) );
AOI22_X1 \dpath/a_mux/_157_ ( .A1(\dpath/a_mux/_063_ ), .A2(\dpath/a_mux/_022_ ), .B1(\dpath/a_mux/_065_ ), .B2(\dpath/a_mux/_038_ ), .ZN(\dpath/a_mux/_060_ ) );
NAND2_X1 \dpath/a_mux/_158_ ( .A1(\dpath/a_mux/_068_ ), .A2(\dpath/a_mux/_006_ ), .ZN(\dpath/a_mux/_061_ ) );
NAND2_X1 \dpath/a_mux/_159_ ( .A1(\dpath/a_mux/_060_ ), .A2(\dpath/a_mux/_061_ ), .ZN(\dpath/a_mux/_093_ ) );
BUF_X1 \dpath/a_mux/_160_ ( .A(\ctrl$a_mux_sel[0] ), .Z(\dpath/a_mux/_103_ ) );
BUF_X1 \dpath/a_mux/_161_ ( .A(\ctrl$a_mux_sel[1] ), .Z(\dpath/a_mux/_104_ ) );
BUF_X1 \dpath/a_mux/_162_ ( .A(\resp_msg[0] ), .Z(\dpath/a_mux/_016_ ) );
BUF_X1 \dpath/a_mux/_163_ ( .A(\dpath/a_lt_b$in1[0] ), .Z(\dpath/a_mux/_032_ ) );
BUF_X1 \dpath/a_mux/_164_ ( .A(\req_msg[16] ), .Z(\dpath/a_mux/_000_ ) );
BUF_X1 \dpath/a_mux/_165_ ( .A(\dpath/a_mux/_087_ ), .Z(\dpath/a_mux$out[0] ) );
BUF_X1 \dpath/a_mux/_166_ ( .A(\resp_msg[1] ), .Z(\dpath/a_mux/_023_ ) );
BUF_X1 \dpath/a_mux/_167_ ( .A(\dpath/a_lt_b$in1[1] ), .Z(\dpath/a_mux/_039_ ) );
BUF_X1 \dpath/a_mux/_168_ ( .A(\req_msg[17] ), .Z(\dpath/a_mux/_007_ ) );
BUF_X1 \dpath/a_mux/_169_ ( .A(\dpath/a_mux/_094_ ), .Z(\dpath/a_mux$out[1] ) );
BUF_X1 \dpath/a_mux/_170_ ( .A(\resp_msg[2] ), .Z(\dpath/a_mux/_024_ ) );
BUF_X1 \dpath/a_mux/_171_ ( .A(\dpath/a_lt_b$in1[2] ), .Z(\dpath/a_mux/_040_ ) );
BUF_X1 \dpath/a_mux/_172_ ( .A(\req_msg[18] ), .Z(\dpath/a_mux/_008_ ) );
BUF_X1 \dpath/a_mux/_173_ ( .A(\dpath/a_mux/_095_ ), .Z(\dpath/a_mux$out[2] ) );
BUF_X1 \dpath/a_mux/_174_ ( .A(\resp_msg[3] ), .Z(\dpath/a_mux/_025_ ) );
BUF_X1 \dpath/a_mux/_175_ ( .A(\dpath/a_lt_b$in1[3] ), .Z(\dpath/a_mux/_041_ ) );
BUF_X1 \dpath/a_mux/_176_ ( .A(\req_msg[19] ), .Z(\dpath/a_mux/_009_ ) );
BUF_X1 \dpath/a_mux/_177_ ( .A(\dpath/a_mux/_096_ ), .Z(\dpath/a_mux$out[3] ) );
BUF_X1 \dpath/a_mux/_178_ ( .A(\resp_msg[4] ), .Z(\dpath/a_mux/_026_ ) );
BUF_X1 \dpath/a_mux/_179_ ( .A(\dpath/a_lt_b$in1[4] ), .Z(\dpath/a_mux/_042_ ) );
BUF_X1 \dpath/a_mux/_180_ ( .A(\req_msg[20] ), .Z(\dpath/a_mux/_010_ ) );
BUF_X1 \dpath/a_mux/_181_ ( .A(\dpath/a_mux/_097_ ), .Z(\dpath/a_mux$out[4] ) );
BUF_X1 \dpath/a_mux/_182_ ( .A(\resp_msg[5] ), .Z(\dpath/a_mux/_027_ ) );
BUF_X1 \dpath/a_mux/_183_ ( .A(\dpath/a_lt_b$in1[5] ), .Z(\dpath/a_mux/_043_ ) );
BUF_X1 \dpath/a_mux/_184_ ( .A(\req_msg[21] ), .Z(\dpath/a_mux/_011_ ) );
BUF_X1 \dpath/a_mux/_185_ ( .A(\dpath/a_mux/_098_ ), .Z(\dpath/a_mux$out[5] ) );
BUF_X1 \dpath/a_mux/_186_ ( .A(\resp_msg[6] ), .Z(\dpath/a_mux/_028_ ) );
BUF_X1 \dpath/a_mux/_187_ ( .A(\dpath/a_lt_b$in1[6] ), .Z(\dpath/a_mux/_044_ ) );
BUF_X1 \dpath/a_mux/_188_ ( .A(\req_msg[22] ), .Z(\dpath/a_mux/_012_ ) );
BUF_X1 \dpath/a_mux/_189_ ( .A(\dpath/a_mux/_099_ ), .Z(\dpath/a_mux$out[6] ) );
BUF_X1 \dpath/a_mux/_190_ ( .A(\resp_msg[7] ), .Z(\dpath/a_mux/_029_ ) );
BUF_X1 \dpath/a_mux/_191_ ( .A(\dpath/a_lt_b$in1[7] ), .Z(\dpath/a_mux/_045_ ) );
BUF_X1 \dpath/a_mux/_192_ ( .A(\req_msg[23] ), .Z(\dpath/a_mux/_013_ ) );
BUF_X1 \dpath/a_mux/_193_ ( .A(\dpath/a_mux/_100_ ), .Z(\dpath/a_mux$out[7] ) );
BUF_X1 \dpath/a_mux/_194_ ( .A(\resp_msg[8] ), .Z(\dpath/a_mux/_030_ ) );
BUF_X1 \dpath/a_mux/_195_ ( .A(\dpath/a_lt_b$in1[8] ), .Z(\dpath/a_mux/_046_ ) );
BUF_X1 \dpath/a_mux/_196_ ( .A(\req_msg[24] ), .Z(\dpath/a_mux/_014_ ) );
BUF_X1 \dpath/a_mux/_197_ ( .A(\dpath/a_mux/_101_ ), .Z(\dpath/a_mux$out[8] ) );
BUF_X1 \dpath/a_mux/_198_ ( .A(\resp_msg[9] ), .Z(\dpath/a_mux/_031_ ) );
BUF_X1 \dpath/a_mux/_199_ ( .A(\dpath/a_lt_b$in1[9] ), .Z(\dpath/a_mux/_047_ ) );
BUF_X1 \dpath/a_mux/_200_ ( .A(\req_msg[25] ), .Z(\dpath/a_mux/_015_ ) );
BUF_X1 \dpath/a_mux/_201_ ( .A(\dpath/a_mux/_102_ ), .Z(\dpath/a_mux$out[9] ) );
BUF_X1 \dpath/a_mux/_202_ ( .A(\resp_msg[10] ), .Z(\dpath/a_mux/_017_ ) );
BUF_X1 \dpath/a_mux/_203_ ( .A(\dpath/a_lt_b$in1[10] ), .Z(\dpath/a_mux/_033_ ) );
BUF_X1 \dpath/a_mux/_204_ ( .A(\req_msg[26] ), .Z(\dpath/a_mux/_001_ ) );
BUF_X1 \dpath/a_mux/_205_ ( .A(\dpath/a_mux/_088_ ), .Z(\dpath/a_mux$out[10] ) );
BUF_X1 \dpath/a_mux/_206_ ( .A(\resp_msg[11] ), .Z(\dpath/a_mux/_018_ ) );
BUF_X1 \dpath/a_mux/_207_ ( .A(\dpath/a_lt_b$in1[11] ), .Z(\dpath/a_mux/_034_ ) );
BUF_X1 \dpath/a_mux/_208_ ( .A(\req_msg[27] ), .Z(\dpath/a_mux/_002_ ) );
BUF_X1 \dpath/a_mux/_209_ ( .A(\dpath/a_mux/_089_ ), .Z(\dpath/a_mux$out[11] ) );
BUF_X1 \dpath/a_mux/_210_ ( .A(\resp_msg[12] ), .Z(\dpath/a_mux/_019_ ) );
BUF_X1 \dpath/a_mux/_211_ ( .A(\dpath/a_lt_b$in1[12] ), .Z(\dpath/a_mux/_035_ ) );
BUF_X1 \dpath/a_mux/_212_ ( .A(\req_msg[28] ), .Z(\dpath/a_mux/_003_ ) );
BUF_X1 \dpath/a_mux/_213_ ( .A(\dpath/a_mux/_090_ ), .Z(\dpath/a_mux$out[12] ) );
BUF_X1 \dpath/a_mux/_214_ ( .A(\resp_msg[13] ), .Z(\dpath/a_mux/_020_ ) );
BUF_X1 \dpath/a_mux/_215_ ( .A(\dpath/a_lt_b$in1[13] ), .Z(\dpath/a_mux/_036_ ) );
BUF_X1 \dpath/a_mux/_216_ ( .A(\req_msg[29] ), .Z(\dpath/a_mux/_004_ ) );
BUF_X1 \dpath/a_mux/_217_ ( .A(\dpath/a_mux/_091_ ), .Z(\dpath/a_mux$out[13] ) );
BUF_X1 \dpath/a_mux/_218_ ( .A(\resp_msg[14] ), .Z(\dpath/a_mux/_021_ ) );
BUF_X1 \dpath/a_mux/_219_ ( .A(\dpath/a_lt_b$in1[14] ), .Z(\dpath/a_mux/_037_ ) );
BUF_X1 \dpath/a_mux/_220_ ( .A(\req_msg[30] ), .Z(\dpath/a_mux/_005_ ) );
BUF_X1 \dpath/a_mux/_221_ ( .A(\dpath/a_mux/_092_ ), .Z(\dpath/a_mux$out[14] ) );
BUF_X1 \dpath/a_mux/_222_ ( .A(\resp_msg[15] ), .Z(\dpath/a_mux/_022_ ) );
BUF_X1 \dpath/a_mux/_223_ ( .A(\dpath/a_lt_b$in1[15] ), .Z(\dpath/a_mux/_038_ ) );
BUF_X1 \dpath/a_mux/_224_ ( .A(\req_msg[31] ), .Z(\dpath/a_mux/_006_ ) );
BUF_X1 \dpath/a_mux/_225_ ( .A(\dpath/a_mux/_093_ ), .Z(\dpath/a_mux$out[15] ) );
MUX2_X1 \dpath/a_reg/_081_ ( .A(\dpath/a_reg/_049_ ), .B(\dpath/a_reg/_033_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_016_ ) );
MUX2_X1 \dpath/a_reg/_082_ ( .A(\dpath/a_reg/_056_ ), .B(\dpath/a_reg/_040_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_023_ ) );
MUX2_X1 \dpath/a_reg/_083_ ( .A(\dpath/a_reg/_057_ ), .B(\dpath/a_reg/_041_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_024_ ) );
MUX2_X1 \dpath/a_reg/_084_ ( .A(\dpath/a_reg/_058_ ), .B(\dpath/a_reg/_042_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_025_ ) );
MUX2_X1 \dpath/a_reg/_085_ ( .A(\dpath/a_reg/_059_ ), .B(\dpath/a_reg/_043_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_026_ ) );
MUX2_X1 \dpath/a_reg/_086_ ( .A(\dpath/a_reg/_060_ ), .B(\dpath/a_reg/_044_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_027_ ) );
MUX2_X1 \dpath/a_reg/_087_ ( .A(\dpath/a_reg/_061_ ), .B(\dpath/a_reg/_045_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_028_ ) );
MUX2_X1 \dpath/a_reg/_088_ ( .A(\dpath/a_reg/_062_ ), .B(\dpath/a_reg/_046_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_029_ ) );
MUX2_X1 \dpath/a_reg/_089_ ( .A(\dpath/a_reg/_063_ ), .B(\dpath/a_reg/_047_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_030_ ) );
MUX2_X1 \dpath/a_reg/_090_ ( .A(\dpath/a_reg/_064_ ), .B(\dpath/a_reg/_048_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_031_ ) );
MUX2_X1 \dpath/a_reg/_091_ ( .A(\dpath/a_reg/_050_ ), .B(\dpath/a_reg/_034_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_017_ ) );
MUX2_X1 \dpath/a_reg/_092_ ( .A(\dpath/a_reg/_051_ ), .B(\dpath/a_reg/_035_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_018_ ) );
MUX2_X1 \dpath/a_reg/_093_ ( .A(\dpath/a_reg/_052_ ), .B(\dpath/a_reg/_036_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_019_ ) );
MUX2_X1 \dpath/a_reg/_094_ ( .A(\dpath/a_reg/_053_ ), .B(\dpath/a_reg/_037_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_020_ ) );
MUX2_X1 \dpath/a_reg/_095_ ( .A(\dpath/a_reg/_054_ ), .B(\dpath/a_reg/_038_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_021_ ) );
MUX2_X1 \dpath/a_reg/_096_ ( .A(\dpath/a_reg/_055_ ), .B(\dpath/a_reg/_039_ ), .S(\dpath/a_reg/_032_ ), .Z(\dpath/a_reg/_022_ ) );
BUF_X1 \dpath/a_reg/_097_ ( .A(\dpath/a_lt_b$in0[0] ), .Z(\dpath/a_reg/_049_ ) );
BUF_X1 \dpath/a_reg/_098_ ( .A(\dpath/a_mux$out[0] ), .Z(\dpath/a_reg/_033_ ) );
BUF_X1 \dpath/a_reg/_099_ ( .A(ctrl$a_reg_en ), .Z(\dpath/a_reg/_032_ ) );
BUF_X1 \dpath/a_reg/_100_ ( .A(\dpath/a_reg/_016_ ), .Z(\dpath/a_reg/_000_ ) );
BUF_X1 \dpath/a_reg/_101_ ( .A(\dpath/a_lt_b$in0[1] ), .Z(\dpath/a_reg/_056_ ) );
BUF_X1 \dpath/a_reg/_102_ ( .A(\dpath/a_mux$out[1] ), .Z(\dpath/a_reg/_040_ ) );
BUF_X1 \dpath/a_reg/_103_ ( .A(\dpath/a_reg/_023_ ), .Z(\dpath/a_reg/_007_ ) );
BUF_X1 \dpath/a_reg/_104_ ( .A(\dpath/a_lt_b$in0[2] ), .Z(\dpath/a_reg/_057_ ) );
BUF_X1 \dpath/a_reg/_105_ ( .A(\dpath/a_mux$out[2] ), .Z(\dpath/a_reg/_041_ ) );
BUF_X1 \dpath/a_reg/_106_ ( .A(\dpath/a_reg/_024_ ), .Z(\dpath/a_reg/_008_ ) );
BUF_X1 \dpath/a_reg/_107_ ( .A(\dpath/a_lt_b$in0[3] ), .Z(\dpath/a_reg/_058_ ) );
BUF_X1 \dpath/a_reg/_108_ ( .A(\dpath/a_mux$out[3] ), .Z(\dpath/a_reg/_042_ ) );
BUF_X1 \dpath/a_reg/_109_ ( .A(\dpath/a_reg/_025_ ), .Z(\dpath/a_reg/_009_ ) );
BUF_X1 \dpath/a_reg/_110_ ( .A(\dpath/a_lt_b$in0[4] ), .Z(\dpath/a_reg/_059_ ) );
BUF_X1 \dpath/a_reg/_111_ ( .A(\dpath/a_mux$out[4] ), .Z(\dpath/a_reg/_043_ ) );
BUF_X1 \dpath/a_reg/_112_ ( .A(\dpath/a_reg/_026_ ), .Z(\dpath/a_reg/_010_ ) );
BUF_X1 \dpath/a_reg/_113_ ( .A(\dpath/a_lt_b$in0[5] ), .Z(\dpath/a_reg/_060_ ) );
BUF_X1 \dpath/a_reg/_114_ ( .A(\dpath/a_mux$out[5] ), .Z(\dpath/a_reg/_044_ ) );
BUF_X1 \dpath/a_reg/_115_ ( .A(\dpath/a_reg/_027_ ), .Z(\dpath/a_reg/_011_ ) );
BUF_X1 \dpath/a_reg/_116_ ( .A(\dpath/a_lt_b$in0[6] ), .Z(\dpath/a_reg/_061_ ) );
BUF_X1 \dpath/a_reg/_117_ ( .A(\dpath/a_mux$out[6] ), .Z(\dpath/a_reg/_045_ ) );
BUF_X1 \dpath/a_reg/_118_ ( .A(\dpath/a_reg/_028_ ), .Z(\dpath/a_reg/_012_ ) );
BUF_X1 \dpath/a_reg/_119_ ( .A(\dpath/a_lt_b$in0[7] ), .Z(\dpath/a_reg/_062_ ) );
BUF_X1 \dpath/a_reg/_120_ ( .A(\dpath/a_mux$out[7] ), .Z(\dpath/a_reg/_046_ ) );
BUF_X1 \dpath/a_reg/_121_ ( .A(\dpath/a_reg/_029_ ), .Z(\dpath/a_reg/_013_ ) );
BUF_X1 \dpath/a_reg/_122_ ( .A(\dpath/a_lt_b$in0[8] ), .Z(\dpath/a_reg/_063_ ) );
BUF_X1 \dpath/a_reg/_123_ ( .A(\dpath/a_mux$out[8] ), .Z(\dpath/a_reg/_047_ ) );
BUF_X1 \dpath/a_reg/_124_ ( .A(\dpath/a_reg/_030_ ), .Z(\dpath/a_reg/_014_ ) );
BUF_X1 \dpath/a_reg/_125_ ( .A(\dpath/a_lt_b$in0[9] ), .Z(\dpath/a_reg/_064_ ) );
BUF_X1 \dpath/a_reg/_126_ ( .A(\dpath/a_mux$out[9] ), .Z(\dpath/a_reg/_048_ ) );
BUF_X1 \dpath/a_reg/_127_ ( .A(\dpath/a_reg/_031_ ), .Z(\dpath/a_reg/_015_ ) );
BUF_X1 \dpath/a_reg/_128_ ( .A(\dpath/a_lt_b$in0[10] ), .Z(\dpath/a_reg/_050_ ) );
BUF_X1 \dpath/a_reg/_129_ ( .A(\dpath/a_mux$out[10] ), .Z(\dpath/a_reg/_034_ ) );
BUF_X1 \dpath/a_reg/_130_ ( .A(\dpath/a_reg/_017_ ), .Z(\dpath/a_reg/_001_ ) );
BUF_X1 \dpath/a_reg/_131_ ( .A(\dpath/a_lt_b$in0[11] ), .Z(\dpath/a_reg/_051_ ) );
BUF_X1 \dpath/a_reg/_132_ ( .A(\dpath/a_mux$out[11] ), .Z(\dpath/a_reg/_035_ ) );
BUF_X1 \dpath/a_reg/_133_ ( .A(\dpath/a_reg/_018_ ), .Z(\dpath/a_reg/_002_ ) );
BUF_X1 \dpath/a_reg/_134_ ( .A(\dpath/a_lt_b$in0[12] ), .Z(\dpath/a_reg/_052_ ) );
BUF_X1 \dpath/a_reg/_135_ ( .A(\dpath/a_mux$out[12] ), .Z(\dpath/a_reg/_036_ ) );
BUF_X1 \dpath/a_reg/_136_ ( .A(\dpath/a_reg/_019_ ), .Z(\dpath/a_reg/_003_ ) );
BUF_X1 \dpath/a_reg/_137_ ( .A(\dpath/a_lt_b$in0[13] ), .Z(\dpath/a_reg/_053_ ) );
BUF_X1 \dpath/a_reg/_138_ ( .A(\dpath/a_mux$out[13] ), .Z(\dpath/a_reg/_037_ ) );
BUF_X1 \dpath/a_reg/_139_ ( .A(\dpath/a_reg/_020_ ), .Z(\dpath/a_reg/_004_ ) );
BUF_X1 \dpath/a_reg/_140_ ( .A(\dpath/a_lt_b$in0[14] ), .Z(\dpath/a_reg/_054_ ) );
BUF_X1 \dpath/a_reg/_141_ ( .A(\dpath/a_mux$out[14] ), .Z(\dpath/a_reg/_038_ ) );
BUF_X1 \dpath/a_reg/_142_ ( .A(\dpath/a_reg/_021_ ), .Z(\dpath/a_reg/_005_ ) );
BUF_X1 \dpath/a_reg/_143_ ( .A(\dpath/a_lt_b$in0[15] ), .Z(\dpath/a_reg/_055_ ) );
BUF_X1 \dpath/a_reg/_144_ ( .A(\dpath/a_mux$out[15] ), .Z(\dpath/a_reg/_039_ ) );
BUF_X1 \dpath/a_reg/_145_ ( .A(\dpath/a_reg/_022_ ), .Z(\dpath/a_reg/_006_ ) );
DFF_X1 \dpath/a_reg/_146_ ( .CK(clk ), .D(\dpath/a_reg/_000_ ), .Q(\dpath/a_lt_b$in0[0] ), .QN(\dpath/a_reg/_065_ ) );
DFF_X1 \dpath/a_reg/_147_ ( .CK(clk ), .D(\dpath/a_reg/_007_ ), .Q(\dpath/a_lt_b$in0[1] ), .QN(\dpath/a_reg/_066_ ) );
DFF_X1 \dpath/a_reg/_148_ ( .CK(clk ), .D(\dpath/a_reg/_008_ ), .Q(\dpath/a_lt_b$in0[2] ), .QN(\dpath/a_reg/_067_ ) );
DFF_X1 \dpath/a_reg/_149_ ( .CK(clk ), .D(\dpath/a_reg/_009_ ), .Q(\dpath/a_lt_b$in0[3] ), .QN(\dpath/a_reg/_068_ ) );
DFF_X1 \dpath/a_reg/_150_ ( .CK(clk ), .D(\dpath/a_reg/_010_ ), .Q(\dpath/a_lt_b$in0[4] ), .QN(\dpath/a_reg/_069_ ) );
DFF_X1 \dpath/a_reg/_151_ ( .CK(clk ), .D(\dpath/a_reg/_011_ ), .Q(\dpath/a_lt_b$in0[5] ), .QN(\dpath/a_reg/_070_ ) );
DFF_X1 \dpath/a_reg/_152_ ( .CK(clk ), .D(\dpath/a_reg/_012_ ), .Q(\dpath/a_lt_b$in0[6] ), .QN(\dpath/a_reg/_071_ ) );
DFF_X1 \dpath/a_reg/_153_ ( .CK(clk ), .D(\dpath/a_reg/_013_ ), .Q(\dpath/a_lt_b$in0[7] ), .QN(\dpath/a_reg/_072_ ) );
DFF_X1 \dpath/a_reg/_154_ ( .CK(clk ), .D(\dpath/a_reg/_014_ ), .Q(\dpath/a_lt_b$in0[8] ), .QN(\dpath/a_reg/_073_ ) );
DFF_X1 \dpath/a_reg/_155_ ( .CK(clk ), .D(\dpath/a_reg/_015_ ), .Q(\dpath/a_lt_b$in0[9] ), .QN(\dpath/a_reg/_074_ ) );
DFF_X1 \dpath/a_reg/_156_ ( .CK(clk ), .D(\dpath/a_reg/_001_ ), .Q(\dpath/a_lt_b$in0[10] ), .QN(\dpath/a_reg/_075_ ) );
DFF_X1 \dpath/a_reg/_157_ ( .CK(clk ), .D(\dpath/a_reg/_002_ ), .Q(\dpath/a_lt_b$in0[11] ), .QN(\dpath/a_reg/_076_ ) );
DFF_X1 \dpath/a_reg/_158_ ( .CK(clk ), .D(\dpath/a_reg/_003_ ), .Q(\dpath/a_lt_b$in0[12] ), .QN(\dpath/a_reg/_077_ ) );
DFF_X1 \dpath/a_reg/_159_ ( .CK(clk ), .D(\dpath/a_reg/_004_ ), .Q(\dpath/a_lt_b$in0[13] ), .QN(\dpath/a_reg/_078_ ) );
DFF_X1 \dpath/a_reg/_160_ ( .CK(clk ), .D(\dpath/a_reg/_005_ ), .Q(\dpath/a_lt_b$in0[14] ), .QN(\dpath/a_reg/_079_ ) );
DFF_X1 \dpath/a_reg/_161_ ( .CK(clk ), .D(\dpath/a_reg/_006_ ), .Q(\dpath/a_lt_b$in0[15] ), .QN(\dpath/a_reg/_080_ ) );
MUX2_X1 \dpath/b_mux/_049_ ( .A(\dpath/b_mux/_000_ ), .B(\dpath/b_mux/_016_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_032_ ) );
MUX2_X1 \dpath/b_mux/_050_ ( .A(\dpath/b_mux/_007_ ), .B(\dpath/b_mux/_023_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_039_ ) );
MUX2_X1 \dpath/b_mux/_051_ ( .A(\dpath/b_mux/_008_ ), .B(\dpath/b_mux/_024_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_040_ ) );
MUX2_X1 \dpath/b_mux/_052_ ( .A(\dpath/b_mux/_009_ ), .B(\dpath/b_mux/_025_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_041_ ) );
MUX2_X1 \dpath/b_mux/_053_ ( .A(\dpath/b_mux/_010_ ), .B(\dpath/b_mux/_026_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_042_ ) );
MUX2_X1 \dpath/b_mux/_054_ ( .A(\dpath/b_mux/_011_ ), .B(\dpath/b_mux/_027_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_043_ ) );
MUX2_X1 \dpath/b_mux/_055_ ( .A(\dpath/b_mux/_012_ ), .B(\dpath/b_mux/_028_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_044_ ) );
MUX2_X1 \dpath/b_mux/_056_ ( .A(\dpath/b_mux/_013_ ), .B(\dpath/b_mux/_029_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_045_ ) );
MUX2_X1 \dpath/b_mux/_057_ ( .A(\dpath/b_mux/_014_ ), .B(\dpath/b_mux/_030_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_046_ ) );
MUX2_X1 \dpath/b_mux/_058_ ( .A(\dpath/b_mux/_015_ ), .B(\dpath/b_mux/_031_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_047_ ) );
MUX2_X1 \dpath/b_mux/_059_ ( .A(\dpath/b_mux/_001_ ), .B(\dpath/b_mux/_017_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_033_ ) );
MUX2_X1 \dpath/b_mux/_060_ ( .A(\dpath/b_mux/_002_ ), .B(\dpath/b_mux/_018_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_034_ ) );
MUX2_X1 \dpath/b_mux/_061_ ( .A(\dpath/b_mux/_003_ ), .B(\dpath/b_mux/_019_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_035_ ) );
MUX2_X1 \dpath/b_mux/_062_ ( .A(\dpath/b_mux/_004_ ), .B(\dpath/b_mux/_020_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_036_ ) );
MUX2_X1 \dpath/b_mux/_063_ ( .A(\dpath/b_mux/_005_ ), .B(\dpath/b_mux/_021_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_037_ ) );
MUX2_X1 \dpath/b_mux/_064_ ( .A(\dpath/b_mux/_006_ ), .B(\dpath/b_mux/_022_ ), .S(\dpath/b_mux/_048_ ), .Z(\dpath/b_mux/_038_ ) );
BUF_X1 \dpath/b_mux/_065_ ( .A(\dpath/a_lt_b$in0[0] ), .Z(\dpath/b_mux/_000_ ) );
BUF_X1 \dpath/b_mux/_066_ ( .A(\req_msg[0] ), .Z(\dpath/b_mux/_016_ ) );
BUF_X1 \dpath/b_mux/_067_ ( .A(ctrl$b_mux_sel ), .Z(\dpath/b_mux/_048_ ) );
BUF_X1 \dpath/b_mux/_068_ ( .A(\dpath/b_mux/_032_ ), .Z(\dpath/b_mux$out[0] ) );
BUF_X1 \dpath/b_mux/_069_ ( .A(\dpath/a_lt_b$in0[1] ), .Z(\dpath/b_mux/_007_ ) );
BUF_X1 \dpath/b_mux/_070_ ( .A(\req_msg[1] ), .Z(\dpath/b_mux/_023_ ) );
BUF_X1 \dpath/b_mux/_071_ ( .A(\dpath/b_mux/_039_ ), .Z(\dpath/b_mux$out[1] ) );
BUF_X1 \dpath/b_mux/_072_ ( .A(\dpath/a_lt_b$in0[2] ), .Z(\dpath/b_mux/_008_ ) );
BUF_X1 \dpath/b_mux/_073_ ( .A(\req_msg[2] ), .Z(\dpath/b_mux/_024_ ) );
BUF_X1 \dpath/b_mux/_074_ ( .A(\dpath/b_mux/_040_ ), .Z(\dpath/b_mux$out[2] ) );
BUF_X1 \dpath/b_mux/_075_ ( .A(\dpath/a_lt_b$in0[3] ), .Z(\dpath/b_mux/_009_ ) );
BUF_X1 \dpath/b_mux/_076_ ( .A(\req_msg[3] ), .Z(\dpath/b_mux/_025_ ) );
BUF_X1 \dpath/b_mux/_077_ ( .A(\dpath/b_mux/_041_ ), .Z(\dpath/b_mux$out[3] ) );
BUF_X1 \dpath/b_mux/_078_ ( .A(\dpath/a_lt_b$in0[4] ), .Z(\dpath/b_mux/_010_ ) );
BUF_X1 \dpath/b_mux/_079_ ( .A(\req_msg[4] ), .Z(\dpath/b_mux/_026_ ) );
BUF_X1 \dpath/b_mux/_080_ ( .A(\dpath/b_mux/_042_ ), .Z(\dpath/b_mux$out[4] ) );
BUF_X1 \dpath/b_mux/_081_ ( .A(\dpath/a_lt_b$in0[5] ), .Z(\dpath/b_mux/_011_ ) );
BUF_X1 \dpath/b_mux/_082_ ( .A(\req_msg[5] ), .Z(\dpath/b_mux/_027_ ) );
BUF_X1 \dpath/b_mux/_083_ ( .A(\dpath/b_mux/_043_ ), .Z(\dpath/b_mux$out[5] ) );
BUF_X1 \dpath/b_mux/_084_ ( .A(\dpath/a_lt_b$in0[6] ), .Z(\dpath/b_mux/_012_ ) );
BUF_X1 \dpath/b_mux/_085_ ( .A(\req_msg[6] ), .Z(\dpath/b_mux/_028_ ) );
BUF_X1 \dpath/b_mux/_086_ ( .A(\dpath/b_mux/_044_ ), .Z(\dpath/b_mux$out[6] ) );
BUF_X1 \dpath/b_mux/_087_ ( .A(\dpath/a_lt_b$in0[7] ), .Z(\dpath/b_mux/_013_ ) );
BUF_X1 \dpath/b_mux/_088_ ( .A(\req_msg[7] ), .Z(\dpath/b_mux/_029_ ) );
BUF_X1 \dpath/b_mux/_089_ ( .A(\dpath/b_mux/_045_ ), .Z(\dpath/b_mux$out[7] ) );
BUF_X1 \dpath/b_mux/_090_ ( .A(\dpath/a_lt_b$in0[8] ), .Z(\dpath/b_mux/_014_ ) );
BUF_X1 \dpath/b_mux/_091_ ( .A(\req_msg[8] ), .Z(\dpath/b_mux/_030_ ) );
BUF_X1 \dpath/b_mux/_092_ ( .A(\dpath/b_mux/_046_ ), .Z(\dpath/b_mux$out[8] ) );
BUF_X1 \dpath/b_mux/_093_ ( .A(\dpath/a_lt_b$in0[9] ), .Z(\dpath/b_mux/_015_ ) );
BUF_X1 \dpath/b_mux/_094_ ( .A(\req_msg[9] ), .Z(\dpath/b_mux/_031_ ) );
BUF_X1 \dpath/b_mux/_095_ ( .A(\dpath/b_mux/_047_ ), .Z(\dpath/b_mux$out[9] ) );
BUF_X1 \dpath/b_mux/_096_ ( .A(\dpath/a_lt_b$in0[10] ), .Z(\dpath/b_mux/_001_ ) );
BUF_X1 \dpath/b_mux/_097_ ( .A(\req_msg[10] ), .Z(\dpath/b_mux/_017_ ) );
BUF_X1 \dpath/b_mux/_098_ ( .A(\dpath/b_mux/_033_ ), .Z(\dpath/b_mux$out[10] ) );
BUF_X1 \dpath/b_mux/_099_ ( .A(\dpath/a_lt_b$in0[11] ), .Z(\dpath/b_mux/_002_ ) );
BUF_X1 \dpath/b_mux/_100_ ( .A(\req_msg[11] ), .Z(\dpath/b_mux/_018_ ) );
BUF_X1 \dpath/b_mux/_101_ ( .A(\dpath/b_mux/_034_ ), .Z(\dpath/b_mux$out[11] ) );
BUF_X1 \dpath/b_mux/_102_ ( .A(\dpath/a_lt_b$in0[12] ), .Z(\dpath/b_mux/_003_ ) );
BUF_X1 \dpath/b_mux/_103_ ( .A(\req_msg[12] ), .Z(\dpath/b_mux/_019_ ) );
BUF_X1 \dpath/b_mux/_104_ ( .A(\dpath/b_mux/_035_ ), .Z(\dpath/b_mux$out[12] ) );
BUF_X1 \dpath/b_mux/_105_ ( .A(\dpath/a_lt_b$in0[13] ), .Z(\dpath/b_mux/_004_ ) );
BUF_X1 \dpath/b_mux/_106_ ( .A(\req_msg[13] ), .Z(\dpath/b_mux/_020_ ) );
BUF_X1 \dpath/b_mux/_107_ ( .A(\dpath/b_mux/_036_ ), .Z(\dpath/b_mux$out[13] ) );
BUF_X1 \dpath/b_mux/_108_ ( .A(\dpath/a_lt_b$in0[14] ), .Z(\dpath/b_mux/_005_ ) );
BUF_X1 \dpath/b_mux/_109_ ( .A(\req_msg[14] ), .Z(\dpath/b_mux/_021_ ) );
BUF_X1 \dpath/b_mux/_110_ ( .A(\dpath/b_mux/_037_ ), .Z(\dpath/b_mux$out[14] ) );
BUF_X1 \dpath/b_mux/_111_ ( .A(\dpath/a_lt_b$in0[15] ), .Z(\dpath/b_mux/_006_ ) );
BUF_X1 \dpath/b_mux/_112_ ( .A(\req_msg[15] ), .Z(\dpath/b_mux/_022_ ) );
BUF_X1 \dpath/b_mux/_113_ ( .A(\dpath/b_mux/_038_ ), .Z(\dpath/b_mux$out[15] ) );
MUX2_X1 \dpath/b_reg/_081_ ( .A(\dpath/b_reg/_049_ ), .B(\dpath/b_reg/_033_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_016_ ) );
MUX2_X1 \dpath/b_reg/_082_ ( .A(\dpath/b_reg/_056_ ), .B(\dpath/b_reg/_040_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_023_ ) );
MUX2_X1 \dpath/b_reg/_083_ ( .A(\dpath/b_reg/_057_ ), .B(\dpath/b_reg/_041_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_024_ ) );
MUX2_X1 \dpath/b_reg/_084_ ( .A(\dpath/b_reg/_058_ ), .B(\dpath/b_reg/_042_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_025_ ) );
MUX2_X1 \dpath/b_reg/_085_ ( .A(\dpath/b_reg/_059_ ), .B(\dpath/b_reg/_043_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_026_ ) );
MUX2_X1 \dpath/b_reg/_086_ ( .A(\dpath/b_reg/_060_ ), .B(\dpath/b_reg/_044_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_027_ ) );
MUX2_X1 \dpath/b_reg/_087_ ( .A(\dpath/b_reg/_061_ ), .B(\dpath/b_reg/_045_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_028_ ) );
MUX2_X1 \dpath/b_reg/_088_ ( .A(\dpath/b_reg/_062_ ), .B(\dpath/b_reg/_046_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_029_ ) );
MUX2_X1 \dpath/b_reg/_089_ ( .A(\dpath/b_reg/_063_ ), .B(\dpath/b_reg/_047_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_030_ ) );
MUX2_X1 \dpath/b_reg/_090_ ( .A(\dpath/b_reg/_064_ ), .B(\dpath/b_reg/_048_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_031_ ) );
MUX2_X1 \dpath/b_reg/_091_ ( .A(\dpath/b_reg/_050_ ), .B(\dpath/b_reg/_034_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_017_ ) );
MUX2_X1 \dpath/b_reg/_092_ ( .A(\dpath/b_reg/_051_ ), .B(\dpath/b_reg/_035_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_018_ ) );
MUX2_X1 \dpath/b_reg/_093_ ( .A(\dpath/b_reg/_052_ ), .B(\dpath/b_reg/_036_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_019_ ) );
MUX2_X1 \dpath/b_reg/_094_ ( .A(\dpath/b_reg/_053_ ), .B(\dpath/b_reg/_037_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_020_ ) );
MUX2_X1 \dpath/b_reg/_095_ ( .A(\dpath/b_reg/_054_ ), .B(\dpath/b_reg/_038_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_021_ ) );
MUX2_X1 \dpath/b_reg/_096_ ( .A(\dpath/b_reg/_055_ ), .B(\dpath/b_reg/_039_ ), .S(\dpath/b_reg/_032_ ), .Z(\dpath/b_reg/_022_ ) );
BUF_X1 \dpath/b_reg/_097_ ( .A(\dpath/a_lt_b$in1[0] ), .Z(\dpath/b_reg/_049_ ) );
BUF_X1 \dpath/b_reg/_098_ ( .A(\dpath/b_mux$out[0] ), .Z(\dpath/b_reg/_033_ ) );
BUF_X1 \dpath/b_reg/_099_ ( .A(ctrl$b_reg_en ), .Z(\dpath/b_reg/_032_ ) );
BUF_X1 \dpath/b_reg/_100_ ( .A(\dpath/b_reg/_016_ ), .Z(\dpath/b_reg/_000_ ) );
BUF_X1 \dpath/b_reg/_101_ ( .A(\dpath/a_lt_b$in1[1] ), .Z(\dpath/b_reg/_056_ ) );
BUF_X1 \dpath/b_reg/_102_ ( .A(\dpath/b_mux$out[1] ), .Z(\dpath/b_reg/_040_ ) );
BUF_X1 \dpath/b_reg/_103_ ( .A(\dpath/b_reg/_023_ ), .Z(\dpath/b_reg/_007_ ) );
BUF_X1 \dpath/b_reg/_104_ ( .A(\dpath/a_lt_b$in1[2] ), .Z(\dpath/b_reg/_057_ ) );
BUF_X1 \dpath/b_reg/_105_ ( .A(\dpath/b_mux$out[2] ), .Z(\dpath/b_reg/_041_ ) );
BUF_X1 \dpath/b_reg/_106_ ( .A(\dpath/b_reg/_024_ ), .Z(\dpath/b_reg/_008_ ) );
BUF_X1 \dpath/b_reg/_107_ ( .A(\dpath/a_lt_b$in1[3] ), .Z(\dpath/b_reg/_058_ ) );
BUF_X1 \dpath/b_reg/_108_ ( .A(\dpath/b_mux$out[3] ), .Z(\dpath/b_reg/_042_ ) );
BUF_X1 \dpath/b_reg/_109_ ( .A(\dpath/b_reg/_025_ ), .Z(\dpath/b_reg/_009_ ) );
BUF_X1 \dpath/b_reg/_110_ ( .A(\dpath/a_lt_b$in1[4] ), .Z(\dpath/b_reg/_059_ ) );
BUF_X1 \dpath/b_reg/_111_ ( .A(\dpath/b_mux$out[4] ), .Z(\dpath/b_reg/_043_ ) );
BUF_X1 \dpath/b_reg/_112_ ( .A(\dpath/b_reg/_026_ ), .Z(\dpath/b_reg/_010_ ) );
BUF_X1 \dpath/b_reg/_113_ ( .A(\dpath/a_lt_b$in1[5] ), .Z(\dpath/b_reg/_060_ ) );
BUF_X1 \dpath/b_reg/_114_ ( .A(\dpath/b_mux$out[5] ), .Z(\dpath/b_reg/_044_ ) );
BUF_X1 \dpath/b_reg/_115_ ( .A(\dpath/b_reg/_027_ ), .Z(\dpath/b_reg/_011_ ) );
BUF_X1 \dpath/b_reg/_116_ ( .A(\dpath/a_lt_b$in1[6] ), .Z(\dpath/b_reg/_061_ ) );
BUF_X1 \dpath/b_reg/_117_ ( .A(\dpath/b_mux$out[6] ), .Z(\dpath/b_reg/_045_ ) );
BUF_X1 \dpath/b_reg/_118_ ( .A(\dpath/b_reg/_028_ ), .Z(\dpath/b_reg/_012_ ) );
BUF_X1 \dpath/b_reg/_119_ ( .A(\dpath/a_lt_b$in1[7] ), .Z(\dpath/b_reg/_062_ ) );
BUF_X1 \dpath/b_reg/_120_ ( .A(\dpath/b_mux$out[7] ), .Z(\dpath/b_reg/_046_ ) );
BUF_X1 \dpath/b_reg/_121_ ( .A(\dpath/b_reg/_029_ ), .Z(\dpath/b_reg/_013_ ) );
BUF_X1 \dpath/b_reg/_122_ ( .A(\dpath/a_lt_b$in1[8] ), .Z(\dpath/b_reg/_063_ ) );
BUF_X1 \dpath/b_reg/_123_ ( .A(\dpath/b_mux$out[8] ), .Z(\dpath/b_reg/_047_ ) );
BUF_X1 \dpath/b_reg/_124_ ( .A(\dpath/b_reg/_030_ ), .Z(\dpath/b_reg/_014_ ) );
BUF_X1 \dpath/b_reg/_125_ ( .A(\dpath/a_lt_b$in1[9] ), .Z(\dpath/b_reg/_064_ ) );
BUF_X1 \dpath/b_reg/_126_ ( .A(\dpath/b_mux$out[9] ), .Z(\dpath/b_reg/_048_ ) );
BUF_X1 \dpath/b_reg/_127_ ( .A(\dpath/b_reg/_031_ ), .Z(\dpath/b_reg/_015_ ) );
BUF_X1 \dpath/b_reg/_128_ ( .A(\dpath/a_lt_b$in1[10] ), .Z(\dpath/b_reg/_050_ ) );
BUF_X1 \dpath/b_reg/_129_ ( .A(\dpath/b_mux$out[10] ), .Z(\dpath/b_reg/_034_ ) );
BUF_X1 \dpath/b_reg/_130_ ( .A(\dpath/b_reg/_017_ ), .Z(\dpath/b_reg/_001_ ) );
BUF_X1 \dpath/b_reg/_131_ ( .A(\dpath/a_lt_b$in1[11] ), .Z(\dpath/b_reg/_051_ ) );
BUF_X1 \dpath/b_reg/_132_ ( .A(\dpath/b_mux$out[11] ), .Z(\dpath/b_reg/_035_ ) );
BUF_X1 \dpath/b_reg/_133_ ( .A(\dpath/b_reg/_018_ ), .Z(\dpath/b_reg/_002_ ) );
BUF_X1 \dpath/b_reg/_134_ ( .A(\dpath/a_lt_b$in1[12] ), .Z(\dpath/b_reg/_052_ ) );
BUF_X1 \dpath/b_reg/_135_ ( .A(\dpath/b_mux$out[12] ), .Z(\dpath/b_reg/_036_ ) );
BUF_X1 \dpath/b_reg/_136_ ( .A(\dpath/b_reg/_019_ ), .Z(\dpath/b_reg/_003_ ) );
BUF_X1 \dpath/b_reg/_137_ ( .A(\dpath/a_lt_b$in1[13] ), .Z(\dpath/b_reg/_053_ ) );
BUF_X1 \dpath/b_reg/_138_ ( .A(\dpath/b_mux$out[13] ), .Z(\dpath/b_reg/_037_ ) );
BUF_X1 \dpath/b_reg/_139_ ( .A(\dpath/b_reg/_020_ ), .Z(\dpath/b_reg/_004_ ) );
BUF_X1 \dpath/b_reg/_140_ ( .A(\dpath/a_lt_b$in1[14] ), .Z(\dpath/b_reg/_054_ ) );
BUF_X1 \dpath/b_reg/_141_ ( .A(\dpath/b_mux$out[14] ), .Z(\dpath/b_reg/_038_ ) );
BUF_X1 \dpath/b_reg/_142_ ( .A(\dpath/b_reg/_021_ ), .Z(\dpath/b_reg/_005_ ) );
BUF_X1 \dpath/b_reg/_143_ ( .A(\dpath/a_lt_b$in1[15] ), .Z(\dpath/b_reg/_055_ ) );
BUF_X1 \dpath/b_reg/_144_ ( .A(\dpath/b_mux$out[15] ), .Z(\dpath/b_reg/_039_ ) );
BUF_X1 \dpath/b_reg/_145_ ( .A(\dpath/b_reg/_022_ ), .Z(\dpath/b_reg/_006_ ) );
DFF_X1 \dpath/b_reg/_146_ ( .CK(clk ), .D(\dpath/b_reg/_000_ ), .Q(\dpath/a_lt_b$in1[0] ), .QN(\dpath/b_reg/_065_ ) );
DFF_X1 \dpath/b_reg/_147_ ( .CK(clk ), .D(\dpath/b_reg/_007_ ), .Q(\dpath/a_lt_b$in1[1] ), .QN(\dpath/b_reg/_066_ ) );
DFF_X1 \dpath/b_reg/_148_ ( .CK(clk ), .D(\dpath/b_reg/_008_ ), .Q(\dpath/a_lt_b$in1[2] ), .QN(\dpath/b_reg/_067_ ) );
DFF_X1 \dpath/b_reg/_149_ ( .CK(clk ), .D(\dpath/b_reg/_009_ ), .Q(\dpath/a_lt_b$in1[3] ), .QN(\dpath/b_reg/_068_ ) );
DFF_X1 \dpath/b_reg/_150_ ( .CK(clk ), .D(\dpath/b_reg/_010_ ), .Q(\dpath/a_lt_b$in1[4] ), .QN(\dpath/b_reg/_069_ ) );
DFF_X1 \dpath/b_reg/_151_ ( .CK(clk ), .D(\dpath/b_reg/_011_ ), .Q(\dpath/a_lt_b$in1[5] ), .QN(\dpath/b_reg/_070_ ) );
DFF_X1 \dpath/b_reg/_152_ ( .CK(clk ), .D(\dpath/b_reg/_012_ ), .Q(\dpath/a_lt_b$in1[6] ), .QN(\dpath/b_reg/_071_ ) );
DFF_X1 \dpath/b_reg/_153_ ( .CK(clk ), .D(\dpath/b_reg/_013_ ), .Q(\dpath/a_lt_b$in1[7] ), .QN(\dpath/b_reg/_072_ ) );
DFF_X1 \dpath/b_reg/_154_ ( .CK(clk ), .D(\dpath/b_reg/_014_ ), .Q(\dpath/a_lt_b$in1[8] ), .QN(\dpath/b_reg/_073_ ) );
DFF_X1 \dpath/b_reg/_155_ ( .CK(clk ), .D(\dpath/b_reg/_015_ ), .Q(\dpath/a_lt_b$in1[9] ), .QN(\dpath/b_reg/_074_ ) );
DFF_X1 \dpath/b_reg/_156_ ( .CK(clk ), .D(\dpath/b_reg/_001_ ), .Q(\dpath/a_lt_b$in1[10] ), .QN(\dpath/b_reg/_075_ ) );
DFF_X1 \dpath/b_reg/_157_ ( .CK(clk ), .D(\dpath/b_reg/_002_ ), .Q(\dpath/a_lt_b$in1[11] ), .QN(\dpath/b_reg/_076_ ) );
DFF_X1 \dpath/b_reg/_158_ ( .CK(clk ), .D(\dpath/b_reg/_003_ ), .Q(\dpath/a_lt_b$in1[12] ), .QN(\dpath/b_reg/_077_ ) );
DFF_X1 \dpath/b_reg/_159_ ( .CK(clk ), .D(\dpath/b_reg/_004_ ), .Q(\dpath/a_lt_b$in1[13] ), .QN(\dpath/b_reg/_078_ ) );
DFF_X1 \dpath/b_reg/_160_ ( .CK(clk ), .D(\dpath/b_reg/_005_ ), .Q(\dpath/a_lt_b$in1[14] ), .QN(\dpath/b_reg/_079_ ) );
DFF_X1 \dpath/b_reg/_161_ ( .CK(clk ), .D(\dpath/b_reg/_006_ ), .Q(\dpath/a_lt_b$in1[15] ), .QN(\dpath/b_reg/_080_ ) );
NOR4_X2 \dpath/b_zero/_21_ ( .A1(\dpath/b_zero/_07_ ), .A2(\dpath/b_zero/_08_ ), .A3(\dpath/b_zero/_10_ ), .A4(\dpath/b_zero/_13_ ), .ZN(\dpath/b_zero/_16_ ) );
NOR4_X2 \dpath/b_zero/_22_ ( .A1(\dpath/b_zero/_14_ ), .A2(\dpath/b_zero/_02_ ), .A3(\dpath/b_zero/_04_ ), .A4(\dpath/b_zero/_05_ ), .ZN(\dpath/b_zero/_17_ ) );
NOR4_X2 \dpath/b_zero/_23_ ( .A1(\dpath/b_zero/_00_ ), .A2(\dpath/b_zero/_09_ ), .A3(\dpath/b_zero/_11_ ), .A4(\dpath/b_zero/_12_ ), .ZN(\dpath/b_zero/_18_ ) );
NOR4_X4 \dpath/b_zero/_24_ ( .A1(\dpath/b_zero/_15_ ), .A2(\dpath/b_zero/_01_ ), .A3(\dpath/b_zero/_03_ ), .A4(\dpath/b_zero/_06_ ), .ZN(\dpath/b_zero/_19_ ) );
AND4_X1 \dpath/b_zero/_25_ ( .A1(\dpath/b_zero/_16_ ), .A2(\dpath/b_zero/_17_ ), .A3(\dpath/b_zero/_18_ ), .A4(\dpath/b_zero/_19_ ), .ZN(\dpath/b_zero/_20_ ) );
BUF_X1 \dpath/b_zero/_26_ ( .A(\dpath/a_lt_b$in1[1] ), .Z(\dpath/b_zero/_07_ ) );
BUF_X1 \dpath/b_zero/_27_ ( .A(\dpath/a_lt_b$in1[0] ), .Z(\dpath/b_zero/_00_ ) );
BUF_X1 \dpath/b_zero/_28_ ( .A(\dpath/a_lt_b$in1[3] ), .Z(\dpath/b_zero/_09_ ) );
BUF_X1 \dpath/b_zero/_29_ ( .A(\dpath/a_lt_b$in1[2] ), .Z(\dpath/b_zero/_08_ ) );
BUF_X1 \dpath/b_zero/_30_ ( .A(\dpath/a_lt_b$in1[5] ), .Z(\dpath/b_zero/_11_ ) );
BUF_X1 \dpath/b_zero/_31_ ( .A(\dpath/a_lt_b$in1[4] ), .Z(\dpath/b_zero/_10_ ) );
BUF_X1 \dpath/b_zero/_32_ ( .A(\dpath/a_lt_b$in1[7] ), .Z(\dpath/b_zero/_13_ ) );
BUF_X1 \dpath/b_zero/_33_ ( .A(\dpath/a_lt_b$in1[6] ), .Z(\dpath/b_zero/_12_ ) );
BUF_X1 \dpath/b_zero/_34_ ( .A(\dpath/a_lt_b$in1[9] ), .Z(\dpath/b_zero/_15_ ) );
BUF_X1 \dpath/b_zero/_35_ ( .A(\dpath/a_lt_b$in1[8] ), .Z(\dpath/b_zero/_14_ ) );
BUF_X1 \dpath/b_zero/_36_ ( .A(\dpath/a_lt_b$in1[11] ), .Z(\dpath/b_zero/_02_ ) );
BUF_X1 \dpath/b_zero/_37_ ( .A(\dpath/a_lt_b$in1[10] ), .Z(\dpath/b_zero/_01_ ) );
BUF_X1 \dpath/b_zero/_38_ ( .A(\dpath/a_lt_b$in1[13] ), .Z(\dpath/b_zero/_04_ ) );
BUF_X1 \dpath/b_zero/_39_ ( .A(\dpath/a_lt_b$in1[12] ), .Z(\dpath/b_zero/_03_ ) );
BUF_X1 \dpath/b_zero/_40_ ( .A(\dpath/a_lt_b$in1[15] ), .Z(\dpath/b_zero/_06_ ) );
BUF_X1 \dpath/b_zero/_41_ ( .A(\dpath/a_lt_b$in1[14] ), .Z(\dpath/b_zero/_05_ ) );
BUF_X1 \dpath/b_zero/_42_ ( .A(\dpath/b_zero/_20_ ), .Z(ctrl$is_b_zero ) );
XOR2_X1 \dpath/sub/_140_ ( .A(\dpath/sub/_000_ ), .B(\dpath/sub/_016_ ), .Z(\dpath/sub/_124_ ) );
XNOR2_X2 \dpath/sub/_141_ ( .A(\dpath/sub/_007_ ), .B(\dpath/sub/_023_ ), .ZN(\dpath/sub/_081_ ) );
INV_X16 \dpath/sub/_142_ ( .A(\dpath/sub/_016_ ), .ZN(\dpath/sub/_082_ ) );
OR3_X1 \dpath/sub/_143_ ( .A1(\dpath/sub/_081_ ), .A2(\dpath/sub/_000_ ), .A3(\dpath/sub/_082_ ), .ZN(\dpath/sub/_083_ ) );
OAI21_X1 \dpath/sub/_144_ ( .A(\dpath/sub/_081_ ), .B1(\dpath/sub/_000_ ), .B2(\dpath/sub/_082_ ), .ZN(\dpath/sub/_084_ ) );
AND2_X1 \dpath/sub/_145_ ( .A1(\dpath/sub/_083_ ), .A2(\dpath/sub/_084_ ), .ZN(\dpath/sub/_131_ ) );
INV_X1 \dpath/sub/_146_ ( .A(\dpath/sub/_023_ ), .ZN(\dpath/sub/_085_ ) );
NAND2_X1 \dpath/sub/_147_ ( .A1(\dpath/sub/_085_ ), .A2(\dpath/sub/_007_ ), .ZN(\dpath/sub/_086_ ) );
XNOR2_X2 \dpath/sub/_148_ ( .A(\dpath/sub/_008_ ), .B(\dpath/sub/_024_ ), .ZN(\dpath/sub/_087_ ) );
INV_X1 \dpath/sub/_149_ ( .A(\dpath/sub/_087_ ), .ZN(\dpath/sub/_088_ ) );
AND3_X1 \dpath/sub/_150_ ( .A1(\dpath/sub/_084_ ), .A2(\dpath/sub/_086_ ), .A3(\dpath/sub/_088_ ), .ZN(\dpath/sub/_089_ ) );
AOI21_X1 \dpath/sub/_151_ ( .A(\dpath/sub/_088_ ), .B1(\dpath/sub/_084_ ), .B2(\dpath/sub/_086_ ), .ZN(\dpath/sub/_090_ ) );
NOR2_X1 \dpath/sub/_152_ ( .A1(\dpath/sub/_089_ ), .A2(\dpath/sub/_090_ ), .ZN(\dpath/sub/_132_ ) );
INV_X1 \dpath/sub/_153_ ( .A(\dpath/sub/_008_ ), .ZN(\dpath/sub/_091_ ) );
NOR2_X2 \dpath/sub/_154_ ( .A1(\dpath/sub/_091_ ), .A2(\dpath/sub/_024_ ), .ZN(\dpath/sub/_092_ ) );
NOR2_X1 \dpath/sub/_155_ ( .A1(\dpath/sub/_090_ ), .A2(\dpath/sub/_092_ ), .ZN(\dpath/sub/_093_ ) );
XNOR2_X2 \dpath/sub/_156_ ( .A(\dpath/sub/_009_ ), .B(\dpath/sub/_025_ ), .ZN(\dpath/sub/_094_ ) );
XNOR2_X1 \dpath/sub/_157_ ( .A(\dpath/sub/_093_ ), .B(\dpath/sub/_094_ ), .ZN(\dpath/sub/_133_ ) );
AND2_X2 \dpath/sub/_158_ ( .A1(\dpath/sub/_094_ ), .A2(\dpath/sub/_092_ ), .ZN(\dpath/sub/_095_ ) );
INV_X1 \dpath/sub/_159_ ( .A(\dpath/sub/_025_ ), .ZN(\dpath/sub/_096_ ) );
AOI21_X4 \dpath/sub/_160_ ( .A(\dpath/sub/_095_ ), .B1(\dpath/sub/_009_ ), .B2(\dpath/sub/_096_ ), .ZN(\dpath/sub/_097_ ) );
INV_X2 \dpath/sub/_161_ ( .A(\dpath/sub/_097_ ), .ZN(\dpath/sub/_098_ ) );
NAND2_X1 \dpath/sub/_162_ ( .A1(\dpath/sub/_087_ ), .A2(\dpath/sub/_094_ ), .ZN(\dpath/sub/_099_ ) );
AOI21_X4 \dpath/sub/_163_ ( .A(\dpath/sub/_099_ ), .B1(\dpath/sub/_084_ ), .B2(\dpath/sub/_086_ ), .ZN(\dpath/sub/_100_ ) );
NOR2_X4 \dpath/sub/_164_ ( .A1(\dpath/sub/_098_ ), .A2(\dpath/sub/_100_ ), .ZN(\dpath/sub/_101_ ) );
XNOR2_X2 \dpath/sub/_165_ ( .A(\dpath/sub/_010_ ), .B(\dpath/sub/_026_ ), .ZN(\dpath/sub/_102_ ) );
XNOR2_X1 \dpath/sub/_166_ ( .A(\dpath/sub/_101_ ), .B(\dpath/sub/_102_ ), .ZN(\dpath/sub/_134_ ) );
INV_X32 \dpath/sub/_167_ ( .A(\dpath/sub/_010_ ), .ZN(\dpath/sub/_103_ ) );
AND2_X1 \dpath/sub/_168_ ( .A1(\dpath/sub/_103_ ), .A2(\dpath/sub/_026_ ), .ZN(\dpath/sub/_104_ ) );
NOR2_X1 \dpath/sub/_169_ ( .A1(\dpath/sub/_103_ ), .A2(\dpath/sub/_026_ ), .ZN(\dpath/sub/_105_ ) );
NOR3_X1 \dpath/sub/_170_ ( .A1(\dpath/sub/_101_ ), .A2(\dpath/sub/_104_ ), .A3(\dpath/sub/_105_ ), .ZN(\dpath/sub/_106_ ) );
NOR2_X1 \dpath/sub/_171_ ( .A1(\dpath/sub/_106_ ), .A2(\dpath/sub/_105_ ), .ZN(\dpath/sub/_107_ ) );
XNOR2_X2 \dpath/sub/_172_ ( .A(\dpath/sub/_011_ ), .B(\dpath/sub/_027_ ), .ZN(\dpath/sub/_108_ ) );
XNOR2_X1 \dpath/sub/_173_ ( .A(\dpath/sub/_107_ ), .B(\dpath/sub/_108_ ), .ZN(\dpath/sub/_135_ ) );
AND2_X1 \dpath/sub/_174_ ( .A1(\dpath/sub/_102_ ), .A2(\dpath/sub/_108_ ), .ZN(\dpath/sub/_109_ ) );
INV_X8 \dpath/sub/_175_ ( .A(\dpath/sub/_109_ ), .ZN(\dpath/sub/_110_ ) );
NOR2_X1 \dpath/sub/_176_ ( .A1(\dpath/sub/_101_ ), .A2(\dpath/sub/_110_ ), .ZN(\dpath/sub/_111_ ) );
INV_X1 \dpath/sub/_177_ ( .A(\dpath/sub/_011_ ), .ZN(\dpath/sub/_112_ ) );
NOR2_X1 \dpath/sub/_178_ ( .A1(\dpath/sub/_112_ ), .A2(\dpath/sub/_027_ ), .ZN(\dpath/sub/_113_ ) );
AOI21_X1 \dpath/sub/_179_ ( .A(\dpath/sub/_113_ ), .B1(\dpath/sub/_108_ ), .B2(\dpath/sub/_105_ ), .ZN(\dpath/sub/_114_ ) );
INV_X1 \dpath/sub/_180_ ( .A(\dpath/sub/_114_ ), .ZN(\dpath/sub/_115_ ) );
XNOR2_X2 \dpath/sub/_181_ ( .A(\dpath/sub/_012_ ), .B(\dpath/sub/_028_ ), .ZN(\dpath/sub/_116_ ) );
OR3_X1 \dpath/sub/_182_ ( .A1(\dpath/sub/_111_ ), .A2(\dpath/sub/_115_ ), .A3(\dpath/sub/_116_ ), .ZN(\dpath/sub/_117_ ) );
OAI21_X1 \dpath/sub/_183_ ( .A(\dpath/sub/_116_ ), .B1(\dpath/sub/_111_ ), .B2(\dpath/sub/_115_ ), .ZN(\dpath/sub/_118_ ) );
AND2_X1 \dpath/sub/_184_ ( .A1(\dpath/sub/_117_ ), .A2(\dpath/sub/_118_ ), .ZN(\dpath/sub/_136_ ) );
INV_X1 \dpath/sub/_185_ ( .A(\dpath/sub/_028_ ), .ZN(\dpath/sub/_119_ ) );
NAND2_X1 \dpath/sub/_186_ ( .A1(\dpath/sub/_119_ ), .A2(\dpath/sub/_012_ ), .ZN(\dpath/sub/_120_ ) );
AND2_X1 \dpath/sub/_187_ ( .A1(\dpath/sub/_118_ ), .A2(\dpath/sub/_120_ ), .ZN(\dpath/sub/_121_ ) );
XNOR2_X2 \dpath/sub/_188_ ( .A(\dpath/sub/_013_ ), .B(\dpath/sub/_029_ ), .ZN(\dpath/sub/_122_ ) );
XNOR2_X1 \dpath/sub/_189_ ( .A(\dpath/sub/_121_ ), .B(\dpath/sub/_122_ ), .ZN(\dpath/sub/_137_ ) );
NAND2_X2 \dpath/sub/_190_ ( .A1(\dpath/sub/_116_ ), .A2(\dpath/sub/_122_ ), .ZN(\dpath/sub/_123_ ) );
NOR3_X4 \dpath/sub/_191_ ( .A1(\dpath/sub/_101_ ), .A2(\dpath/sub/_110_ ), .A3(\dpath/sub/_123_ ), .ZN(\dpath/sub/_032_ ) );
NAND3_X1 \dpath/sub/_192_ ( .A1(\dpath/sub/_122_ ), .A2(\dpath/sub/_012_ ), .A3(\dpath/sub/_119_ ), .ZN(\dpath/sub/_033_ ) );
INV_X1 \dpath/sub/_193_ ( .A(\dpath/sub/_013_ ), .ZN(\dpath/sub/_034_ ) );
OAI221_X4 \dpath/sub/_194_ ( .A(\dpath/sub/_033_ ), .B1(\dpath/sub/_034_ ), .B2(\dpath/sub/_029_ ), .C1(\dpath/sub/_114_ ), .C2(\dpath/sub/_123_ ), .ZN(\dpath/sub/_035_ ) );
NOR2_X4 \dpath/sub/_195_ ( .A1(\dpath/sub/_032_ ), .A2(\dpath/sub/_035_ ), .ZN(\dpath/sub/_036_ ) );
XNOR2_X2 \dpath/sub/_196_ ( .A(\dpath/sub/_014_ ), .B(\dpath/sub/_030_ ), .ZN(\dpath/sub/_037_ ) );
XNOR2_X1 \dpath/sub/_197_ ( .A(\dpath/sub/_036_ ), .B(\dpath/sub/_037_ ), .ZN(\dpath/sub/_138_ ) );
OAI21_X1 \dpath/sub/_198_ ( .A(\dpath/sub/_037_ ), .B1(\dpath/sub/_032_ ), .B2(\dpath/sub/_035_ ), .ZN(\dpath/sub/_038_ ) );
INV_X1 \dpath/sub/_199_ ( .A(\dpath/sub/_014_ ), .ZN(\dpath/sub/_039_ ) );
NOR2_X2 \dpath/sub/_200_ ( .A1(\dpath/sub/_039_ ), .A2(\dpath/sub/_030_ ), .ZN(\dpath/sub/_040_ ) );
INV_X1 \dpath/sub/_201_ ( .A(\dpath/sub/_040_ ), .ZN(\dpath/sub/_041_ ) );
AND2_X1 \dpath/sub/_202_ ( .A1(\dpath/sub/_038_ ), .A2(\dpath/sub/_041_ ), .ZN(\dpath/sub/_042_ ) );
XNOR2_X2 \dpath/sub/_203_ ( .A(\dpath/sub/_015_ ), .B(\dpath/sub/_031_ ), .ZN(\dpath/sub/_043_ ) );
XNOR2_X1 \dpath/sub/_204_ ( .A(\dpath/sub/_042_ ), .B(\dpath/sub/_043_ ), .ZN(\dpath/sub/_139_ ) );
OAI211_X2 \dpath/sub/_205_ ( .A(\dpath/sub/_037_ ), .B(\dpath/sub/_043_ ), .C1(\dpath/sub/_032_ ), .C2(\dpath/sub/_035_ ), .ZN(\dpath/sub/_044_ ) );
AND2_X2 \dpath/sub/_206_ ( .A1(\dpath/sub/_043_ ), .A2(\dpath/sub/_040_ ), .ZN(\dpath/sub/_045_ ) );
INV_X1 \dpath/sub/_207_ ( .A(\dpath/sub/_031_ ), .ZN(\dpath/sub/_046_ ) );
AOI21_X4 \dpath/sub/_208_ ( .A(\dpath/sub/_045_ ), .B1(\dpath/sub/_015_ ), .B2(\dpath/sub/_046_ ), .ZN(\dpath/sub/_047_ ) );
AND2_X2 \dpath/sub/_209_ ( .A1(\dpath/sub/_044_ ), .A2(\dpath/sub/_047_ ), .ZN(\dpath/sub/_048_ ) );
XNOR2_X1 \dpath/sub/_210_ ( .A(\dpath/sub/_001_ ), .B(\dpath/sub/_017_ ), .ZN(\dpath/sub/_049_ ) );
XNOR2_X1 \dpath/sub/_211_ ( .A(\dpath/sub/_048_ ), .B(\dpath/sub/_049_ ), .ZN(\dpath/sub/_125_ ) );
INV_X1 \dpath/sub/_212_ ( .A(\dpath/sub/_001_ ), .ZN(\dpath/sub/_050_ ) );
NOR2_X1 \dpath/sub/_213_ ( .A1(\dpath/sub/_050_ ), .A2(\dpath/sub/_017_ ), .ZN(\dpath/sub/_051_ ) );
AND2_X1 \dpath/sub/_214_ ( .A1(\dpath/sub/_050_ ), .A2(\dpath/sub/_017_ ), .ZN(\dpath/sub/_052_ ) );
NOR3_X2 \dpath/sub/_215_ ( .A1(\dpath/sub/_048_ ), .A2(\dpath/sub/_051_ ), .A3(\dpath/sub/_052_ ), .ZN(\dpath/sub/_053_ ) );
NOR2_X2 \dpath/sub/_216_ ( .A1(\dpath/sub/_053_ ), .A2(\dpath/sub/_051_ ), .ZN(\dpath/sub/_054_ ) );
XNOR2_X1 \dpath/sub/_217_ ( .A(\dpath/sub/_002_ ), .B(\dpath/sub/_018_ ), .ZN(\dpath/sub/_055_ ) );
XNOR2_X1 \dpath/sub/_218_ ( .A(\dpath/sub/_054_ ), .B(\dpath/sub/_055_ ), .ZN(\dpath/sub/_126_ ) );
NAND4_X1 \dpath/sub/_219_ ( .A1(\dpath/sub/_037_ ), .A2(\dpath/sub/_043_ ), .A3(\dpath/sub/_049_ ), .A4(\dpath/sub/_055_ ), .ZN(\dpath/sub/_056_ ) );
NOR2_X4 \dpath/sub/_220_ ( .A1(\dpath/sub/_036_ ), .A2(\dpath/sub/_056_ ), .ZN(\dpath/sub/_057_ ) );
NAND2_X1 \dpath/sub/_221_ ( .A1(\dpath/sub/_055_ ), .A2(\dpath/sub/_051_ ), .ZN(\dpath/sub/_058_ ) );
INV_X1 \dpath/sub/_222_ ( .A(\dpath/sub/_002_ ), .ZN(\dpath/sub/_059_ ) );
NAND2_X1 \dpath/sub/_223_ ( .A1(\dpath/sub/_049_ ), .A2(\dpath/sub/_055_ ), .ZN(\dpath/sub/_060_ ) );
OAI221_X4 \dpath/sub/_224_ ( .A(\dpath/sub/_058_ ), .B1(\dpath/sub/_059_ ), .B2(\dpath/sub/_018_ ), .C1(\dpath/sub/_047_ ), .C2(\dpath/sub/_060_ ), .ZN(\dpath/sub/_061_ ) );
NOR2_X1 \dpath/sub/_225_ ( .A1(\dpath/sub/_057_ ), .A2(\dpath/sub/_061_ ), .ZN(\dpath/sub/_062_ ) );
XNOR2_X1 \dpath/sub/_226_ ( .A(\dpath/sub/_003_ ), .B(\dpath/sub/_019_ ), .ZN(\dpath/sub/_063_ ) );
XNOR2_X1 \dpath/sub/_227_ ( .A(\dpath/sub/_062_ ), .B(\dpath/sub/_063_ ), .ZN(\dpath/sub/_127_ ) );
OAI21_X1 \dpath/sub/_228_ ( .A(\dpath/sub/_063_ ), .B1(\dpath/sub/_057_ ), .B2(\dpath/sub/_061_ ), .ZN(\dpath/sub/_064_ ) );
INV_X1 \dpath/sub/_229_ ( .A(\dpath/sub/_003_ ), .ZN(\dpath/sub/_065_ ) );
NOR2_X1 \dpath/sub/_230_ ( .A1(\dpath/sub/_065_ ), .A2(\dpath/sub/_019_ ), .ZN(\dpath/sub/_066_ ) );
INV_X1 \dpath/sub/_231_ ( .A(\dpath/sub/_066_ ), .ZN(\dpath/sub/_067_ ) );
AND2_X2 \dpath/sub/_232_ ( .A1(\dpath/sub/_064_ ), .A2(\dpath/sub/_067_ ), .ZN(\dpath/sub/_068_ ) );
XNOR2_X1 \dpath/sub/_233_ ( .A(\dpath/sub/_004_ ), .B(\dpath/sub/_020_ ), .ZN(\dpath/sub/_069_ ) );
XNOR2_X1 \dpath/sub/_234_ ( .A(\dpath/sub/_068_ ), .B(\dpath/sub/_069_ ), .ZN(\dpath/sub/_128_ ) );
OAI211_X4 \dpath/sub/_235_ ( .A(\dpath/sub/_063_ ), .B(\dpath/sub/_069_ ), .C1(\dpath/sub/_057_ ), .C2(\dpath/sub/_061_ ), .ZN(\dpath/sub/_070_ ) );
AND2_X1 \dpath/sub/_236_ ( .A1(\dpath/sub/_069_ ), .A2(\dpath/sub/_066_ ), .ZN(\dpath/sub/_071_ ) );
INV_X1 \dpath/sub/_237_ ( .A(\dpath/sub/_020_ ), .ZN(\dpath/sub/_072_ ) );
AOI21_X1 \dpath/sub/_238_ ( .A(\dpath/sub/_071_ ), .B1(\dpath/sub/_004_ ), .B2(\dpath/sub/_072_ ), .ZN(\dpath/sub/_073_ ) );
XOR2_X1 \dpath/sub/_239_ ( .A(\dpath/sub/_005_ ), .B(\dpath/sub/_021_ ), .Z(\dpath/sub/_074_ ) );
AND3_X1 \dpath/sub/_240_ ( .A1(\dpath/sub/_070_ ), .A2(\dpath/sub/_073_ ), .A3(\dpath/sub/_074_ ), .ZN(\dpath/sub/_075_ ) );
AOI21_X4 \dpath/sub/_241_ ( .A(\dpath/sub/_074_ ), .B1(\dpath/sub/_070_ ), .B2(\dpath/sub/_073_ ), .ZN(\dpath/sub/_076_ ) );
NOR2_X1 \dpath/sub/_242_ ( .A1(\dpath/sub/_075_ ), .A2(\dpath/sub/_076_ ), .ZN(\dpath/sub/_129_ ) );
INV_X1 \dpath/sub/_243_ ( .A(\dpath/sub/_005_ ), .ZN(\dpath/sub/_077_ ) );
NOR2_X1 \dpath/sub/_244_ ( .A1(\dpath/sub/_077_ ), .A2(\dpath/sub/_021_ ), .ZN(\dpath/sub/_078_ ) );
NOR2_X2 \dpath/sub/_245_ ( .A1(\dpath/sub/_076_ ), .A2(\dpath/sub/_078_ ), .ZN(\dpath/sub/_079_ ) );
XNOR2_X1 \dpath/sub/_246_ ( .A(\dpath/sub/_006_ ), .B(\dpath/sub/_022_ ), .ZN(\dpath/sub/_080_ ) );
XNOR2_X1 \dpath/sub/_247_ ( .A(\dpath/sub/_079_ ), .B(\dpath/sub/_080_ ), .ZN(\dpath/sub/_130_ ) );
BUF_X1 \dpath/sub/_248_ ( .A(\dpath/a_lt_b$in0[0] ), .Z(\dpath/sub/_000_ ) );
BUF_X1 \dpath/sub/_249_ ( .A(\dpath/a_lt_b$in1[0] ), .Z(\dpath/sub/_016_ ) );
BUF_X1 \dpath/sub/_250_ ( .A(\dpath/sub/_124_ ), .Z(\resp_msg[0] ) );
BUF_X1 \dpath/sub/_251_ ( .A(\dpath/a_lt_b$in0[1] ), .Z(\dpath/sub/_007_ ) );
BUF_X1 \dpath/sub/_252_ ( .A(\dpath/a_lt_b$in1[1] ), .Z(\dpath/sub/_023_ ) );
BUF_X1 \dpath/sub/_253_ ( .A(\dpath/sub/_131_ ), .Z(\resp_msg[1] ) );
BUF_X1 \dpath/sub/_254_ ( .A(\dpath/a_lt_b$in0[2] ), .Z(\dpath/sub/_008_ ) );
BUF_X1 \dpath/sub/_255_ ( .A(\dpath/a_lt_b$in1[2] ), .Z(\dpath/sub/_024_ ) );
BUF_X1 \dpath/sub/_256_ ( .A(\dpath/sub/_132_ ), .Z(\resp_msg[2] ) );
BUF_X1 \dpath/sub/_257_ ( .A(\dpath/a_lt_b$in0[3] ), .Z(\dpath/sub/_009_ ) );
BUF_X1 \dpath/sub/_258_ ( .A(\dpath/a_lt_b$in1[3] ), .Z(\dpath/sub/_025_ ) );
BUF_X1 \dpath/sub/_259_ ( .A(\dpath/sub/_133_ ), .Z(\resp_msg[3] ) );
BUF_X1 \dpath/sub/_260_ ( .A(\dpath/a_lt_b$in0[4] ), .Z(\dpath/sub/_010_ ) );
BUF_X1 \dpath/sub/_261_ ( .A(\dpath/a_lt_b$in1[4] ), .Z(\dpath/sub/_026_ ) );
BUF_X1 \dpath/sub/_262_ ( .A(\dpath/sub/_134_ ), .Z(\resp_msg[4] ) );
BUF_X1 \dpath/sub/_263_ ( .A(\dpath/a_lt_b$in0[5] ), .Z(\dpath/sub/_011_ ) );
BUF_X1 \dpath/sub/_264_ ( .A(\dpath/a_lt_b$in1[5] ), .Z(\dpath/sub/_027_ ) );
BUF_X1 \dpath/sub/_265_ ( .A(\dpath/sub/_135_ ), .Z(\resp_msg[5] ) );
BUF_X1 \dpath/sub/_266_ ( .A(\dpath/a_lt_b$in0[6] ), .Z(\dpath/sub/_012_ ) );
BUF_X1 \dpath/sub/_267_ ( .A(\dpath/a_lt_b$in1[6] ), .Z(\dpath/sub/_028_ ) );
BUF_X1 \dpath/sub/_268_ ( .A(\dpath/sub/_136_ ), .Z(\resp_msg[6] ) );
BUF_X1 \dpath/sub/_269_ ( .A(\dpath/a_lt_b$in0[7] ), .Z(\dpath/sub/_013_ ) );
BUF_X1 \dpath/sub/_270_ ( .A(\dpath/a_lt_b$in1[7] ), .Z(\dpath/sub/_029_ ) );
BUF_X1 \dpath/sub/_271_ ( .A(\dpath/sub/_137_ ), .Z(\resp_msg[7] ) );
BUF_X1 \dpath/sub/_272_ ( .A(\dpath/a_lt_b$in0[8] ), .Z(\dpath/sub/_014_ ) );
BUF_X1 \dpath/sub/_273_ ( .A(\dpath/a_lt_b$in1[8] ), .Z(\dpath/sub/_030_ ) );
BUF_X1 \dpath/sub/_274_ ( .A(\dpath/sub/_138_ ), .Z(\resp_msg[8] ) );
BUF_X1 \dpath/sub/_275_ ( .A(\dpath/a_lt_b$in0[9] ), .Z(\dpath/sub/_015_ ) );
BUF_X1 \dpath/sub/_276_ ( .A(\dpath/a_lt_b$in1[9] ), .Z(\dpath/sub/_031_ ) );
BUF_X1 \dpath/sub/_277_ ( .A(\dpath/sub/_139_ ), .Z(\resp_msg[9] ) );
BUF_X1 \dpath/sub/_278_ ( .A(\dpath/a_lt_b$in0[10] ), .Z(\dpath/sub/_001_ ) );
BUF_X1 \dpath/sub/_279_ ( .A(\dpath/a_lt_b$in1[10] ), .Z(\dpath/sub/_017_ ) );
BUF_X1 \dpath/sub/_280_ ( .A(\dpath/sub/_125_ ), .Z(\resp_msg[10] ) );
BUF_X1 \dpath/sub/_281_ ( .A(\dpath/a_lt_b$in0[11] ), .Z(\dpath/sub/_002_ ) );
BUF_X1 \dpath/sub/_282_ ( .A(\dpath/a_lt_b$in1[11] ), .Z(\dpath/sub/_018_ ) );
BUF_X1 \dpath/sub/_283_ ( .A(\dpath/sub/_126_ ), .Z(\resp_msg[11] ) );
BUF_X1 \dpath/sub/_284_ ( .A(\dpath/a_lt_b$in0[12] ), .Z(\dpath/sub/_003_ ) );
BUF_X1 \dpath/sub/_285_ ( .A(\dpath/a_lt_b$in1[12] ), .Z(\dpath/sub/_019_ ) );
BUF_X1 \dpath/sub/_286_ ( .A(\dpath/sub/_127_ ), .Z(\resp_msg[12] ) );
BUF_X1 \dpath/sub/_287_ ( .A(\dpath/a_lt_b$in0[13] ), .Z(\dpath/sub/_004_ ) );
BUF_X1 \dpath/sub/_288_ ( .A(\dpath/a_lt_b$in1[13] ), .Z(\dpath/sub/_020_ ) );
BUF_X1 \dpath/sub/_289_ ( .A(\dpath/sub/_128_ ), .Z(\resp_msg[13] ) );
BUF_X1 \dpath/sub/_290_ ( .A(\dpath/a_lt_b$in0[14] ), .Z(\dpath/sub/_005_ ) );
BUF_X1 \dpath/sub/_291_ ( .A(\dpath/a_lt_b$in1[14] ), .Z(\dpath/sub/_021_ ) );
BUF_X1 \dpath/sub/_292_ ( .A(\dpath/sub/_129_ ), .Z(\resp_msg[14] ) );
BUF_X1 \dpath/sub/_293_ ( .A(\dpath/a_lt_b$in0[15] ), .Z(\dpath/sub/_006_ ) );
BUF_X1 \dpath/sub/_294_ ( .A(\dpath/a_lt_b$in1[15] ), .Z(\dpath/sub/_022_ ) );
BUF_X1 \dpath/sub/_295_ ( .A(\dpath/sub/_130_ ), .Z(\resp_msg[15] ) );

endmodule
